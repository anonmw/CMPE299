module dcache_vector(address, data_in, read, write, data_out, valid, CLK, RST);
    parameter WIDTH = 32;
    parameter VEC_WIDTH = 64;
    reg [VEC_WIDTH-1:0] dcache [127:0];
    
    input wire [WIDTH-1:0] address;
    input wire [VEC_WIDTH-1:0] data_in;
    input wire read, write;
    output wire [VEC_WIDTH-1:0] data_out;
    output wire valid;
    input CLK, RST;
    
    assign valid = 1'b1;
    
    wire [6:0] index = address[9:3];
    
    //always do this no matter what (read always active basically)
    assign data_out = dcache[index];
    
    always @ (posedge CLK or posedge RST) begin
        if (RST == 1) begin
            dcache[0] <= 64'h0000000000000000;
            dcache[1] <= 64'h0000000000000001;
            dcache[2] <= 64'h0000000000000002;
            dcache[3] <= 64'h0000000000000003;
            dcache[4] <= 64'h0004000400040004;
            dcache[5] <= 64'h0005000500050005;
            dcache[6] <= 64'h0006000600060006;
            dcache[7] <= 64'h0007000700070007;
            dcache[8] <= 64'h0000000000000008;
            dcache[9] <= 64'h0000000000000009;
            dcache[10] <= 64'h000000000000000A;
            dcache[11] <= 64'h000000000000000B;
            dcache[12] <= 64'h000000000000000C;
            dcache[13] <= 64'h000000000000000D;
            dcache[14] <= 64'h000000000000000E;
            dcache[15] <= 64'h000000000000000F;
            dcache[16] <= 64'h0000000000000000;
            dcache[17] <= 64'h0000000000000000;
            dcache[18] <= 64'h0000000000000000;
            dcache[19] <= 64'h0000000000000000;
            dcache[20] <= 64'h0000000000000000;
            dcache[21] <= 64'h0000000000000000;
            dcache[22] <= 64'h0000000000000000;
            dcache[23] <= 64'h0000000000000000;
            dcache[24] <= 64'h0000000000000000;
            dcache[25] <= 64'h0000000000000000;
            dcache[26] <= 64'h0000000000000000;
            dcache[27] <= 64'h0000000000000000;
            dcache[28] <= 64'h0000000000000000;
            dcache[29] <= 64'h0000000000000000;
            dcache[30] <= 64'h0000000000000000;
            dcache[31] <= 64'h0000000000000000;
            dcache[32] <= 64'h0000000000000000;
            dcache[33] <= 64'h0000000000000001;
            dcache[34] <= 64'h0000000000000002;
            dcache[35] <= 64'h0000000000000003;
            dcache[36] <= 64'h0000000000000004;
            dcache[37] <= 64'h0000000000000005;
            dcache[38] <= 64'h0000000000000006;
            dcache[39] <= 64'h0000000000000007;
            dcache[40] <= 64'h0000000000000008;
            dcache[41] <= 64'h0000000000000009;
            dcache[42] <= 64'h000000000000000A;
            dcache[43] <= 64'h000000000000000B;
            dcache[44] <= 64'h000000000000000C;
            dcache[45] <= 64'h000000000000000D;
            dcache[46] <= 64'h000000000000000E;
            dcache[47] <= 64'h000000000000000F;
            dcache[48] <= 64'h0000000000000000;
            dcache[49] <= 64'h0000000000000000;
            dcache[50] <= 64'h0000000000000000;
            dcache[51] <= 64'h0000000000000000;
            dcache[52] <= 64'h0000000000000000;
            dcache[53] <= 64'h0000000000000000;
            dcache[54] <= 64'h0000000000000000;
            dcache[55] <= 64'h0000000000000000;
            dcache[56] <= 64'h0000000000000000;
            dcache[57] <= 64'h0000000000000000;
            dcache[58] <= 64'h0000000000000000;
            dcache[59] <= 64'h0000000000000000;
            dcache[60] <= 64'h0000000000000000;
            dcache[61] <= 64'h0000000000000000;
            dcache[62] <= 64'h0000000000000000;
            dcache[63] <= 64'h0000000000000000;
            dcache[64] <= 64'h0000000000000000;
            dcache[65] <= 64'h0000000000000001;
            dcache[66] <= 64'h0000000000000002;
            dcache[67] <= 64'h0000000000000003;
            dcache[68] <= 64'h0000000000000004;
            dcache[69] <= 64'h0000000000000005;
            dcache[70] <= 64'h0000000000000006;
            dcache[71] <= 64'h0000000000000007;
            dcache[72] <= 64'h0000000000000008;
            dcache[73] <= 64'h0000000000000009;
            dcache[74] <= 64'h000000000000000A;
            dcache[75] <= 64'h000000000000000B;
            dcache[76] <= 64'h000000000000000C;
            dcache[77] <= 64'h000000000000000D;
            dcache[78] <= 64'h000000000000000E;
            dcache[79] <= 64'h000000000000000F;
            dcache[80] <= 64'h0000000000000000;
            dcache[81] <= 64'h0000000000000000;
            dcache[82] <= 64'h0000000000000000;
            dcache[83] <= 64'h0000000000000000;
            dcache[84] <= 64'h0000000000000000;
            dcache[85] <= 64'h0000000000000000;
            dcache[86] <= 64'h0000000000000000;
            dcache[87] <= 64'h0000000000000000;
            dcache[88] <= 64'h0000000000000000;
            dcache[89] <= 64'h0000000000000000;
            dcache[90] <= 64'h0000000000000000;
            dcache[91] <= 64'h0000000000000000;
            dcache[92] <= 64'h0000000000000000;
            dcache[93] <= 64'h0000000000000000;
            dcache[94] <= 64'h0000000000000000;
            dcache[95] <= 64'h0000000000000000;
            dcache[96] <= 64'h0000000000000000;
            dcache[97] <= 64'h0000000000000001;
            dcache[98] <= 64'h0000000000000002;
            dcache[99] <= 64'h0000000000000003;
            dcache[100] <= 64'h0000000000000004;
            dcache[101] <= 64'h0000000000000005;
            dcache[102] <= 64'h0000000000000006;
            dcache[103] <= 64'h0000000000000007;
            dcache[104] <= 64'h0000000000000008;
            dcache[105] <= 64'h0000000000000009;
            dcache[106] <= 64'h000000000000000A;
            dcache[107] <= 64'h000000000000000B;
            dcache[108] <= 64'h000000000000000C;
            dcache[109] <= 64'h000000000000000D;
            dcache[110] <= 64'h000000000000000E;
            dcache[111] <= 64'h000000000000000F;
            dcache[112] <= 64'h0000000000000000;
            dcache[113] <= 64'h0000000000000000;
            dcache[114] <= 64'h0000000000000000;
            dcache[115] <= 64'h0000000000000000;
            dcache[116] <= 64'h0000000000000000;
            dcache[117] <= 64'h0000000000000000;
            dcache[118] <= 64'h0000000000000000;
            dcache[119] <= 64'h0000000000000000;
            dcache[120] <= 64'h0000000000000000;
            dcache[121] <= 64'h0000000000000000;
            dcache[122] <= 64'h0000000000000000;
            dcache[123] <= 64'h0000000000000000;
            dcache[124] <= 64'h0000000000000000;
            dcache[125] <= 64'h0000000000000000;
            dcache[126] <= 64'h0000000000000000;
            dcache[127] <= 64'h0000000000000000;
        end else if (write == 1) begin
            dcache[index] <= data_in;
        // update value
        end
    end

    initial begin
        $dumpfile("main_tb.vcd");
        $dumpvars(0, dcache[0]);
        $dumpvars(0, dcache[1]);
        $dumpvars(0, dcache[2]);
        $dumpvars(0, dcache[3]);
        $dumpvars(0, dcache[4]);
        $dumpvars(0, dcache[5]);
        $dumpvars(0, dcache[6]);
        $dumpvars(0, dcache[7]);
        $dumpvars(0, dcache[8]);
        $dumpvars(0, dcache[9]);
        $dumpvars(0, dcache[10]);
        $dumpvars(0, dcache[11]);
        $dumpvars(0, dcache[12]);
        $dumpvars(0, dcache[13]);
        $dumpvars(0, dcache[14]);
        $dumpvars(0, dcache[15]);
        $dumpvars(0, dcache[16]);
        $dumpvars(0, dcache[17]);
        $dumpvars(0, dcache[18]);
        $dumpvars(0, dcache[19]);
        $dumpvars(0, dcache[20]);
        $dumpvars(0, dcache[21]);
        $dumpvars(0, dcache[22]);
        $dumpvars(0, dcache[23]);
        $dumpvars(0, dcache[24]);
        $dumpvars(0, dcache[25]);
        $dumpvars(0, dcache[26]);
        $dumpvars(0, dcache[27]);
        $dumpvars(0, dcache[28]);
        $dumpvars(0, dcache[29]);
        $dumpvars(0, dcache[30]);
        $dumpvars(0, dcache[31]);
        $dumpvars(0, dcache[32]);
        $dumpvars(0, dcache[33]);
        $dumpvars(0, dcache[34]);
        $dumpvars(0, dcache[35]);
        $dumpvars(0, dcache[36]);
        $dumpvars(0, dcache[37]);
        $dumpvars(0, dcache[38]);
        $dumpvars(0, dcache[39]);
        $dumpvars(0, dcache[40]);
        $dumpvars(0, dcache[41]);
        $dumpvars(0, dcache[42]);
        $dumpvars(0, dcache[43]);
        $dumpvars(0, dcache[44]);
        $dumpvars(0, dcache[45]);
        $dumpvars(0, dcache[46]);
        $dumpvars(0, dcache[47]);
        $dumpvars(0, dcache[48]);
        $dumpvars(0, dcache[49]);
        $dumpvars(0, dcache[50]);
        $dumpvars(0, dcache[51]);
        $dumpvars(0, dcache[52]);
        $dumpvars(0, dcache[53]);
        $dumpvars(0, dcache[54]);
        $dumpvars(0, dcache[55]);
        $dumpvars(0, dcache[56]);
        $dumpvars(0, dcache[57]);
        $dumpvars(0, dcache[58]);
        $dumpvars(0, dcache[59]);
        $dumpvars(0, dcache[60]);
        $dumpvars(0, dcache[61]);
        $dumpvars(0, dcache[62]);
        $dumpvars(0, dcache[63]);
        $dumpvars(0, dcache[64]);
        $dumpvars(0, dcache[65]);
        $dumpvars(0, dcache[66]);
        $dumpvars(0, dcache[67]);
        $dumpvars(0, dcache[68]);
        $dumpvars(0, dcache[69]);
        $dumpvars(0, dcache[70]);
        $dumpvars(0, dcache[71]);
        $dumpvars(0, dcache[72]);
        $dumpvars(0, dcache[73]);
        $dumpvars(0, dcache[74]);
        $dumpvars(0, dcache[75]);
        $dumpvars(0, dcache[76]);
        $dumpvars(0, dcache[77]);
        $dumpvars(0, dcache[78]);
        $dumpvars(0, dcache[79]);
        $dumpvars(0, dcache[80]);
        $dumpvars(0, dcache[81]);
        $dumpvars(0, dcache[82]);
        $dumpvars(0, dcache[83]);
        $dumpvars(0, dcache[84]);
        $dumpvars(0, dcache[85]);
        $dumpvars(0, dcache[86]);
        $dumpvars(0, dcache[87]);
        $dumpvars(0, dcache[88]);
        $dumpvars(0, dcache[89]);
        $dumpvars(0, dcache[90]);
        $dumpvars(0, dcache[91]);
        $dumpvars(0, dcache[92]);
        $dumpvars(0, dcache[93]);
        $dumpvars(0, dcache[94]);
        $dumpvars(0, dcache[95]);
        $dumpvars(0, dcache[96]);
        $dumpvars(0, dcache[97]);
        $dumpvars(0, dcache[98]);
        $dumpvars(0, dcache[99]);
        $dumpvars(0, dcache[100]);
        $dumpvars(0, dcache[101]);
        $dumpvars(0, dcache[102]);
        $dumpvars(0, dcache[103]);
        $dumpvars(0, dcache[104]);
        $dumpvars(0, dcache[105]);
        $dumpvars(0, dcache[106]);
        $dumpvars(0, dcache[107]);
        $dumpvars(0, dcache[108]);
        $dumpvars(0, dcache[109]);
        $dumpvars(0, dcache[110]);
        $dumpvars(0, dcache[111]);
        $dumpvars(0, dcache[112]);
        $dumpvars(0, dcache[113]);
        $dumpvars(0, dcache[114]);
        $dumpvars(0, dcache[115]);
        $dumpvars(0, dcache[116]);
        $dumpvars(0, dcache[117]);
        $dumpvars(0, dcache[118]);
        $dumpvars(0, dcache[119]);
        $dumpvars(0, dcache[120]);
        $dumpvars(0, dcache[121]);
        $dumpvars(0, dcache[122]);
        $dumpvars(0, dcache[123]);
        $dumpvars(0, dcache[124]);
        $dumpvars(0, dcache[125]);
        $dumpvars(0, dcache[126]);
        $dumpvars(0, dcache[127]);
    end

endmodule
