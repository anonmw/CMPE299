module icache(PC, instruction, CLK, RST);
    parameter WIDTH = 32;
    reg [WIDTH-1:0] icache [127:0];
    
    input wire [WIDTH-1:0] PC;
    output wire [WIDTH-1:0] instruction;
    input wire CLK, RST;
    
    wire [6:0] index = PC[8:2];
    
    assign instruction = icache[index];
    `define TEST_MATMUL
    always @ (posedge CLK or posedge RST) begin
    	if (RST == 1) begin
    	`ifdef TEST_ADDI
    	    icache[0] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1
    	    icache[1] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 2
    	    icache[2] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 3
    	    icache[3] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 4
    	    icache[4] <= 32'b111111111000_00001_000_00001_0010011; // addi r1, r1, -8 #r1 = -4
    	    icache[5] <= 32'b000000010000_00001_000_00001_0010011; // addi r1, r1, 16 #r1 = 12
    	    icache[6] <= 32'b111111110100_00001_000_00001_0010011; // addi r1, r1, -12 #r1 = 0
    	    icache[7] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SLTI
    	    icache[0] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1
    	    icache[1] <= 32'b000000000000_00001_010_00010_0010011; // slti r2, r1, 0 #r2 = 0
    	    icache[2] <= 32'b000000000001_00001_010_00011_0010011; // slti r3, r1, 1 #r3 = 0
    	    icache[3] <= 32'b000000000010_00001_010_00100_0010011; // slti r4, r1, 2 #r4 = 1
    	    icache[4] <= 32'b111111111110_00000_000_00001_0010011; // addi r1, r0, -2 #r1 = -2
    	    icache[5] <= 32'b111111111111_00001_010_00010_0010011; // slti r2, r1, -1 # r2 = 1
    	    icache[6] <= 32'b111111111101_00001_010_00011_0010011; // slti r2, r1, -3 # r3 = 0
    	    icache[7] <= 32'b000000000000_00001_010_00100_0010011; // slti r2, r1, 0 # r4 = 1
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SLTIU
    	    icache[0] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1
    	    icache[1] <= 32'b000000000000_00001_011_00010_0010011; // slti r2, r1, 0 #r2 = 0
    	    icache[2] <= 32'b000000000001_00001_011_00011_0010011; // slti r3, r1, 1 #r3 = 0
    	    icache[3] <= 32'b000000000010_00001_011_00100_0010011; // slti r4, r1, 2 #r4 = 1
    	    icache[4] <= 32'b111111111110_00000_000_00001_0010011; // addi r1, r0, -2 #r1 = -2
    	    icache[5] <= 32'b111111111111_00001_011_00010_0010011; // slti r2, r1, -1 # r2 = 1
    	    icache[6] <= 32'b111111111101_00001_011_00011_0010011; // slti r2, r1, -3 # r3 = 0
    	    icache[7] <= 32'b000000000000_00001_011_00100_0010011; // slti r2, r1, 0 # r4 = 0
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_ANDI
    	    icache[0] <= 32'b010101010101_00000_000_00001_0010011; // addi r1, r0, 1365 #r1 = 1365
    	    icache[1] <= 32'b110101010101_00001_111_00010_0010011; // andi r2, r1, -683 #r2 = 1365
    	    icache[2] <= 32'b010101010101_00001_111_00011_0010011; // andi r3, r1, 1365 #r3 = 1365
    	    icache[3] <= 32'b101010101010_00001_111_00100_0010011; // andi r4, r1, -1366 #r4 = 0
    	    icache[4] <= 32'b101010101010_00000_000_00001_0010011; // addi r1, r0, -1366 #r1 = -1366
    	    icache[5] <= 32'b111111111111_00001_111_00010_0010011; // andi r2, r1, -1 # r2 = -1366
    	    icache[6] <= 32'b001010101010_00001_111_00011_0010011; // andi r2, r1, 682 # r3 = 682
    	    icache[7] <= 32'b010101010101_00001_111_00100_0010011; // andi r2, r1, 341 # r4 = 0
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_ORI
    	    icache[0] <= 32'b010101010101_00000_000_00001_0010011; // addi r1, r0, 1365 #r1 = 1365
    	    icache[1] <= 32'b110101010101_00001_110_00010_0010011; // ori r2, r1, -683 #r2 = -683
    	    icache[2] <= 32'b010101010101_00001_110_00011_0010011; // ori r3, r1, 1365 #r3 = 1365
    	    icache[3] <= 32'b101010101010_00001_110_00100_0010011; // ori r4, r1, -1366 #r4 = -1
    	    icache[4] <= 32'b101010101010_00000_000_00001_0010011; // addi r1, r0, -1366 #r1 = -1366
    	    icache[5] <= 32'b111111111111_00001_110_00010_0010011; // ori r2, r1, -1 # r2 = -1
    	    icache[6] <= 32'b001010101010_00001_110_00011_0010011; // ori r2, r1, 682 # r3 = -1366
    	    icache[7] <= 32'b010101010101_00001_110_00100_0010011; // ori r2, r1, 341 # r4 = -1
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_XORI
    	    icache[0] <= 32'b010101010101_00000_000_00001_0010011; // addi r1, r0, 1365 #r1 = 1365
    	    icache[1] <= 32'b110101010101_00001_100_00010_0010011; // xori r2, r1, -683 #r2 = -2048
    	    icache[2] <= 32'b010101010101_00001_100_00011_0010011; // xori r3, r1, 1365 #r3 = 0
    	    icache[3] <= 32'b101010101010_00001_100_00100_0010011; // xori r4, r1, -1366 #r4 = -1
    	    icache[4] <= 32'b101010101010_00000_000_00001_0010011; // addi r1, r0, -1366 #r1 = -1366
    	    icache[5] <= 32'b111111111111_00001_100_00010_0010011; // xori r2, r1, -1 # r2 = 1365
    	    icache[6] <= 32'b001010101010_00001_100_00011_0010011; // xori r2, r1, 682 # r3 = -2048
    	    icache[7] <= 32'b010101010101_00001_100_00100_0010011; // xori r2, r1, 341 # r4 = -1
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SLLI
    	    icache[0] <= 32'b010101010101_00000_000_00001_0010011; // addi r1, r0, 1365 #r1 = 1365
    	    icache[1] <= 32'b0000000_00001_00001_001_00010_0010011; // slli r2, r1, 1 #r2 = 2730
    	    icache[2] <= 32'b0000000_01000_00001_001_00011_0010011; // slli r3, r1, 8 #r3 = 349440
    	    icache[3] <= 32'b0000000_10000_00001_001_00100_0010011; // slli r4, r1, 16 #r4 = 89456640
    	    icache[4] <= 32'b101010101010_00000_000_00001_0010011; // addi r1, r0, -1366 #r1 = -1366
    	    icache[5] <= 32'b0000000_00001_00001_001_00010_0010011; // slli r2, r1, 1 # r2 = -2732
    	    icache[6] <= 32'b0000000_01000_00001_001_00011_0010011; // slli r2, r1, 8 # r3 = -349696
    	    icache[7] <= 32'b0000000_10000_00001_001_00100_0010011; // slli r2, r1, 16 # r4 = -89522176
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SRLI
    	    icache[0] <= 32'b010101010101_00000_000_00001_0010011; // addi r1, r0, 1365 #r1 = 1365
    	    icache[1] <= 32'b0000000_00001_00001_101_00010_0010011; // srli r2, r1, 1 #r2 = 682
    	    icache[2] <= 32'b0000000_01000_00001_101_00011_0010011; // srli r3, r1, 8 #r3 = 5
    	    icache[3] <= 32'b0000000_10000_00001_101_00100_0010011; // srli r4, r1, 16 #r4 = 0
    	    icache[4] <= 32'b101010101010_00000_000_00001_0010011; // addi r1, r0, -1366 #r1 = -1366
    	    icache[5] <= 32'b0000000_00001_00001_101_00010_0010011; // srli r2, r1, 1 # r2 = 2147482965
    	    icache[6] <= 32'b0000000_01000_00001_101_00011_0010011; // srli r2, r1, 8 # r3 = 16777210
    	    icache[7] <= 32'b0000000_10000_00001_101_00100_0010011; // srli r2, r1, 16 # r4 = 65535
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SRAI
    	    icache[0] <= 32'b010101010101_00000_000_00001_0010011; // addi r1, r0, 1365 #r1 = 1365
    	    icache[1] <= 32'b0100000_00001_00001_101_00010_0010011; // srai r2, r1, 1 #r2 = 682
    	    icache[2] <= 32'b0100000_01000_00001_101_00011_0010011; // srai r3, r1, 8 #r3 = 5
    	    icache[3] <= 32'b0100000_10000_00001_101_00100_0010011; // srai r4, r1, 16 #r4 = 0
    	    icache[4] <= 32'b101010101010_00000_000_00001_0010011; // addi r1, r0, -1366 #r1 = -1366
    	    icache[5] <= 32'b0100000_00001_00001_101_00010_0010011; // srai r2, r1, 1 # r2 = -683
    	    icache[6] <= 32'b0100000_01000_00001_101_00011_0010011; // srai r2, r1, 8 # r3 = -6
    	    icache[7] <= 32'b0100000_10000_00001_101_00100_0010011; // srai r2, r1, 16 # r4 = -1
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_LUI_AUIPC
    	    icache[0] <= 32'b01010101010100000000_00001_0110111; // lui r1, 349696 #r1 = 1431306240
    	    icache[1] <= 32'b11111111111111111111_00010_0110111; // lui r2, -1 #r2 = -4096
    	    icache[2] <= 32'b10000000000000000000_00011_0110111; // lui r3, -524288 #r3 = -2147483648
    	    icache[3] <= 32'b00000000000000000000_00100_0110111; // lui r4, 0 #r4 = 0
    	    icache[4] <= 32'b00000000000000000000_00101_0010111; // auipc r5, 0 #r1 = 16
    	    icache[5] <= 32'b11111111111111111111_00110_0010111; // auipc r6, 1 # r2 = -4076
    	    icache[6] <= 32'b10000000000000000000_00111_0010111; // auipc r7, -524288 # r3 = -2147483624
    	    icache[7] <= 32'b00000000000000000001_01000_0010111; // auipc r8, 1 # r4 = 4124
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_ADD
    	    icache[0] <= 32'b000000000010_00000_000_00001_0010011; // addi r1, r0, 2 #r1 = 2
    	    icache[1] <= 32'b000000000011_00000_000_00010_0010011; // addi r2, r0, 3 #r2 = 3
    	    icache[2] <= 32'b111111111110_00000_000_00011_0010011; // addi r3, r0, -2 #r3 = -2
    	    icache[3] <= 32'b111111111101_00000_000_00100_0010011; // addi r4, r0, -3 #r4 = -3
    	    icache[4] <= 32'b0000000_00010_00001_000_00101_0110011; // add r5, r1, r2 #r5 = 5
    	    icache[5] <= 32'b0000000_00100_00001_000_00110_0110011; // add r6, r1, r4 #r6 = -1
    	    icache[6] <= 32'b0000000_00011_00010_000_00111_0110011; // add r7, r2, r3 #r7 = 1
    	    icache[7] <= 32'b0000000_00100_00011_000_01000_0110011; // add r8, r3, r4 #r8 = -5
    	    icache[8] <= 32'b0000000_00001_00011_000_01001_0110011; // add r9, r3, r1 #r9 = 0
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SUB
    	    icache[0] <= 32'b000000000010_00000_000_00001_0010011; // addi r1, r0, 2 #r1 = 2
    	    icache[1] <= 32'b000000000011_00000_000_00010_0010011; // addi r2, r0, 3 #r2 = 3
    	    icache[2] <= 32'b111111111110_00000_000_00011_0010011; // addi r3, r0, -2 #r3 = -2
    	    icache[3] <= 32'b111111111101_00000_000_00100_0010011; // addi r4, r0, -3 #r4 = -3
    	    icache[4] <= 32'b0100000_00010_00001_000_00101_0110011; // sub r5, r1, r2 #r5 = 2-3= -1
    	    icache[5] <= 32'b0100000_00001_00010_000_00110_0110011; // sub r6, r2, r1 #r6 = 3-2= 1
    	    icache[6] <= 32'b0100000_00100_00011_000_00111_0110011; // sub r7, r3, r4 #r7 = -2-(-)3 = 1
    	    icache[7] <= 32'b0100000_00011_00100_000_01000_0110011; // sub r8, r4, r3 #r8 = -3-(-2) = -1
    	    icache[8] <= 32'b0100000_00011_00001_000_01001_0110011; // sub r9, r1, r3 #r9 = 2-(-2)= 4
    	    icache[9] <= 32'b0100000_00001_00011_000_01010_0110011; // sub r10, r3, r1 #r10 = -2-2= -4
    	    icache[10] <= 32'b0100000_00001_00001_000_01011_0110011; // sub r11, r1, r1 #r11 = 2-2 = 0
    	    icache[11] <= 32'b0100000_00011_00011_000_01100_0110011; // sub r12, r3, r3 #r12 = -2-(-2) = 0
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SLT
    	    icache[0] <= 32'b000000000010_00000_000_00001_0010011; // addi r1, r0, 2 #r1 = 2
    	    icache[1] <= 32'b000000000011_00000_000_00010_0010011; // addi r2, r0, 3 #r2 = 3
    	    icache[2] <= 32'b111111111110_00000_000_00011_0010011; // addi r3, r0, -2 #r3 = -2
    	    icache[3] <= 32'b111111111101_00000_000_00100_0010011; // addi r4, r0, -3 #r4 = -3
    	    icache[4] <= 32'b0000000_00010_00001_010_00101_0110011; // slt r5, r1, r2 #r5 = 2<3=1
    	    icache[5] <= 32'b0000000_00001_00010_010_00110_0110011; // slt r6, r2, r1 #r6 = 3<2=0
    	    icache[6] <= 32'b0000000_00001_00001_010_00111_0110011; // slt r7, r1, r1 #r7 = 2<2=0
    	    icache[7] <= 32'b0000000_00011_00001_010_01000_0110011; // slt r8, r1, r3 #r8 = 2<-2=0
    	    icache[8] <= 32'b0000000_00100_00001_010_01001_0110011; // slt r9, r1, r4 #r9 = 2<-3= 0
    	    icache[9] <= 32'b0000000_00001_00011_010_01010_0110011; // slt r10, r3, r1 #r10 = -2<2= 1
    	    icache[10] <= 32'b0000000_00010_00011_010_01011_0110011; // slt r11, r3, r2 #r11 = -2<3 = 1
    	    icache[11] <= 32'b0000000_00011_00100_010_01100_0110011; // slt r12, r4, r3 #r12 = -3<-2 = 1
    	    icache[12] <= 32'b0000000_00100_00011_010_01101_0110011; // slt r13, r3, r4 #r13 = -2<-3 = 0
    	    icache[13] <= 32'b0000000_00011_00011_010_01110_0110011; // slt r14, r3, r3 #r14 = -2<-2 = 0
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SLTU
    	    icache[0] <= 32'b000000000010_00000_000_00001_0010011; // addi r1, r0, 2 #r1 = 2
    	    icache[1] <= 32'b000000000011_00000_000_00010_0010011; // addi r2, r0, 3 #r2 = 3
    	    icache[2] <= 32'b111111111110_00000_000_00011_0010011; // addi r3, r0, -2 #r3 = -2
    	    icache[3] <= 32'b111111111101_00000_000_00100_0010011; // addi r4, r0, -3 #r4 = -3
    	    icache[4] <= 32'b0100000_00010_00001_011_00101_0110011; // sltu r5, r1, r2 #r5 = 2<3=1
    	    icache[5] <= 32'b0100000_00001_00010_011_00110_0110011; // sltu r6, r2, r1 #r6 = 3<2=0
    	    icache[6] <= 32'b0100000_00001_00001_011_00111_0110011; // sltu r7, r1, r1 #r7 = 2<2=0
    	    icache[7] <= 32'b0100000_00011_00001_011_01000_0110011; // sltu r8, r1, r3 #r8 = 2<-2=1
    	    icache[8] <= 32'b0100000_00100_00001_011_01001_0110011; // sltu r9, r1, r4 #r9 = 2<-3= 1
    	    icache[9] <= 32'b0100000_00001_00011_011_01010_0110011; // sltu r10, r3, r1 #r10 = -2<2= 0
    	    icache[10] <= 32'b0100000_00010_00011_011_01011_0110011; // sltu r11, r3, r2 #r11 = -2<3 = 0
    	    icache[11] <= 32'b0100000_00011_00100_011_01100_0110011; // sltu r12, r4, r3 #r12 = -3<-2 = 1
    	    icache[12] <= 32'b0100000_00100_00011_011_01101_0110011; // sltu r13, r3, r4 #r13 = -2<-3 = 0
    	    icache[13] <= 32'b0100000_00011_00011_011_01110_0110011; // sltu r14, r3, r3 #r14 = -2<-2 = 0
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_AND
    	    icache[0] <= 32'b01010101010101010101_00001_0110111; // lui r1, 0x55555 #r1 = 0x55555000
    	    icache[1] <= 32'b010101010101_00001_000_00001_0010011; // addi r1, r1, 0x555 #r1 = 0x55555555
    	    icache[2] <= 32'b10101010101010101010_00010_0110111; // lui r2, 0xAAAAA #r1 = 0xAAAAA000
    	    icache[3] <= 32'b010000000000_00010_000_00010_0010011; // addi r2, r2, 0x400 #r2 = 0xAAAAA400
    	    icache[4] <= 32'b011010101010_00010_000_00010_0010011; // addi r2, r2, 0x6AA #r2 = 0xAAAAAAAA
    	    icache[5] <= 32'b111111111111_00000_000_00011_0010011; // addi r3, r0, -1 #r3 = 0xFFFFFFFF
    	    icache[6] <= 32'b0000000_00010_00001_111_00100_0110011; // and r4, r1, r2 #r4 = 0
    	    icache[7] <= 32'b0000000_00001_00001_111_00101_0110011; // and r5, r1, r1 #r5 = 0x55555555
    	    icache[8] <= 32'b0000000_00011_00001_111_00110_0110011; // and r6, r1, r3 #r6 = 0x55555555
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_OR
    	    icache[0] <= 32'b01010101010101010101_00001_0110111; // lui r1, 0x55555 #r1 = 0x55555000
    	    icache[1] <= 32'b010101010101_00001_000_00001_0010011; // addi r1, r1, 0x555 #r1 = 0x55555555
    	    icache[2] <= 32'b10101010101010101010_00010_0110111; // lui r2, 0xAAAAA #r1 = 0xAAAAA000
    	    icache[3] <= 32'b010000000000_00010_000_00010_0010011; // addi r2, r2, 0x400 #r2 = 0xAAAAA400
    	    icache[4] <= 32'b011010101010_00010_000_00010_0010011; // addi r2, r2, 0x6AA #r2 = 0xAAAAAAAA
    	    icache[5] <= 32'b111111111111_00000_000_00011_0010011; // addi r3, r0, -1 #r3 = 0xFFFFFFFF
    	    icache[6] <= 32'b0000000_00010_00001_110_00100_0110011; // or r4, r1, r2 #r4 = 0xFFFFFFFF
    	    icache[7] <= 32'b0000000_00001_00001_110_00101_0110011; // or r5, r1, r1 #r5 = 0x55555555
    	    icache[8] <= 32'b0000000_00011_00001_110_00110_0110011; // or r6, r1, r3 #r6 = 0xFFFFFFFF
    	    icache[9] <= 32'b0000000_00000_00001_110_00111_0110011; // or r7, r1, r0 #r7 = 0x55555555
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_XOR
    	    icache[0] <= 32'b01010101010101010101_00001_0110111; // lui r1, 0x55555 #r1 = 0x55555000
    	    icache[1] <= 32'b010101010101_00001_000_00001_0010011; // addi r1, r1, 0x555 #r1 = 0x55555555
    	    icache[2] <= 32'b10101010101010101010_00010_0110111; // lui r2, 0xAAAAA #r1 = 0xAAAAA000
    	    icache[3] <= 32'b010000000000_00010_000_00010_0010011; // addi r2, r2, 0x400 #r2 = 0xAAAAA400
    	    icache[4] <= 32'b011010101010_00010_000_00010_0010011; // addi r2, r2, 0x6AA #r2 = 0xAAAAAAAA
    	    icache[5] <= 32'b111111111111_00000_000_00011_0010011; // addi r3, r0, -1 #r3 = 0xFFFFFFFF
    	    icache[6] <= 32'b0000000_00010_00001_100_00100_0110011; // xor r4, r1, r2 #r4 = 0xFFFFFFFF
    	    icache[7] <= 32'b0000000_00001_00001_100_00101_0110011; // xor r5, r1, r1 #r5 = 0x00000000
    	    icache[8] <= 32'b0000000_00011_00001_100_00110_0110011; // xor r6, r1, r3 #r6 = 0xAAAAAAAA
    	    icache[9] <= 32'b0000000_00000_00001_100_00111_0110011; // xor r7, r1, r0 #r7 = 0x55555555
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SLL
    	    icache[0] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1
    	    icache[1] <= 32'b000000001000_00000_000_00010_0010011; // addi r2, r0, 8 #r2 = 8
    	    icache[2] <= 32'b000000010000_00000_000_00011_0010011; // addi r3, r0, 16 #r3 = 16
    	    icache[3] <= 32'b111111111111_00000_000_00100_0010011; // addi r4, r0, -1 #r4 = 0xFFFFFFFF
    	    icache[4] <= 32'b0000000_00001_00100_001_00101_0110011; // sll r5, r4, r1 #r5 = 0xFFFFFFFE
    	    icache[5] <= 32'b0000000_00010_00100_001_00110_0110011; // sll r6, r4, r2 #r6 = 0xFFFFFF00
    	    icache[6] <= 32'b0000000_00011_00100_001_00111_0110011; // sll r7, r4, r3 #r7 = 0xFFFF0000
    	    icache[7] <= 32'b0000000_00011_00111_001_01000_0110011; // sll r8, r7, r3 #r8 = 0x00000000
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SRL
    	    icache[0] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1
    	    icache[1] <= 32'b000000001000_00000_000_00010_0010011; // addi r2, r0, 8 #r2 = 8
    	    icache[2] <= 32'b000000010000_00000_000_00011_0010011; // addi r3, r0, 16 #r3 = 16
    	    icache[3] <= 32'b111111111111_00000_000_00100_0010011; // addi r4, r0, -1 #r4 = 0xFFFFFFFF
    	    icache[4] <= 32'b0000000_00001_00100_101_00101_0110011; // srl r5, r4, r1 #r5 = 0x7FFFFFFF
    	    icache[5] <= 32'b0000000_00010_00100_101_00110_0110011; // srl r6, r4, r2 #r6 = 0x00FFFFFF
    	    icache[6] <= 32'b0000000_00011_00100_101_00111_0110011; // srl r7, r4, r3 #r7 = 0x0000FFFF
    	    icache[7] <= 32'b0000000_00011_00111_101_01000_0110011; // srl r8, r7, r3 #r8 = 0x00000000
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_SRA
    	    icache[0] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1
    	    icache[1] <= 32'b000000001000_00000_000_00010_0010011; // addi r2, r0, 8 #r2 = 8
    	    icache[2] <= 32'b000000010000_00000_000_00011_0010011; // addi r3, r0, 16 #r3 = 16
    	    icache[3] <= 32'b111111111111_00000_000_00100_0010011; // addi r4, r0, -1 #r4 = 0xFFFFFFFF
    	    icache[4] <= 32'b0100000_00001_00100_101_00101_0110011; // srl r5, r4, r1 #r5 = 0xFFFFFFFF
    	    icache[5] <= 32'b0100000_00010_00100_101_00110_0110011; // srl r6, r4, r2 #r6 = 0xFFFFFFFF
    	    icache[6] <= 32'b0100000_00011_00100_101_00111_0110011; // srl r7, r4, r3 #r7 = 0xFFFFFFFF
    	    icache[7] <= 32'b0100000_00011_00111_101_01000_0110011; // srl r8, r7, r3 #r8 = 0xFFFFFFFF
    	    icache[8] <= 32'b10000000000000000000_01001_0110111; // lui r9, 0x80000 #r9 = 0x80000000
    	    icache[9] <= 32'b0100000_00001_01001_101_01010_0110011; // srl r10, r9, r1 #r10 = 0xC0000000
    	    icache[10] <= 32'b0100000_00010_01001_101_01011_0110011; // srl r11, r9, r2 #r11 = 0xFF800000
    	    icache[11] <= 32'b0100000_00011_01001_101_01100_0110011; // srl r12, r9, r3 #r12 = 0xFFFF8000
    	    icache[12] <= 32'b0100000_00011_01100_101_01101_0110011; // srl r13, r12, r3 #r13 = 0xFFFFFFFF
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
	    `endif
    	`ifdef TEST_JAL
    	    icache[0] <= 32'b000000000000_00000_000_00001_0010011; // addi r1, r0, 0 #r1 = 0
    	    icache[1] <= 32'b0_0000000100_0_00000000_00010_1101111; // jal r2, 8 #r2 = 8
    	    icache[2] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1 # shouldn't happen, jumped over
    	    icache[3] <= 32'b0_0000000100_0_00000000_00011_1101111; // jal r3, 8 #r3 = 16
    	    icache[4] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1 # shouldn't happen, jumped over
    	    icache[5] <= 32'b0_0000000100_0_00000000_00100_1101111; // jal r4, 8 #r4 = 24
    	    icache[6] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1 # shouldn't happen, jumped over
    	    icache[7] <= 32'b0_0000000110_0_00000000_00101_1101111; // jal r5, 12 #r5 = 32
    	    icache[8] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1 # shouldn't happen, jumped over
    	    icache[9] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1 # shouldn't happen, jumped over
    	    icache[10] <= 32'b0_0000001010_0_00000000_00110_1101111; // jal r6, 20 #r6 = 44
    	    icache[11] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r0, 1 #r1 = 1 # r1 = 1
    	    icache[12] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r0, 1 #r1 = 1 # r1 = 2
    	    icache[13] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r0, 1 #r1 = 1 # r1 = 3
    	    icache[14] <= 32'b1_1111100100_1_11111111_01000_1101111; // jal r8, -56 #r8 = 60
    	    icache[15] <= 32'b1_1111111000_1_11111111_00111_1101111; // jal r7, -16 #r7 = 64
	    `endif
    	`ifdef TEST_JALR
    	    icache[0] <= 32'b000000101000_00000_000_00001_0010011; // addi r1, r0, 40 #r1 = 40
    	    icache[1] <= 32'b000000001100_00000_000_00010_1100111; // jalr r2, r0, 12 #r2 = 8
    	    icache[2] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # shouldn't happen, jumped over
    	    icache[3] <= 32'b111111101100_00001_000_00011_1100111; // jalr r3, r1, -20 #r3 = 16
    	    icache[4] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # shouldn't happen, jumped over
    	    icache[5] <= 32'b111111110100_00001_000_00100_1100111; // jalr r4, r1, -12 #r4 = 24
    	    icache[6] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # shouldn't happen, jumped over
    	    icache[7] <= 32'b000000000000_00001_000_00101_1100111; // jalr r5, r0, 0 #r5 = 32
    	    icache[8] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # shouldn't happen, jumped over
    	    icache[9] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # shouldn't happen, jumped over
    	    icache[10] <= 32'b00000010100_00001_000_00010_1100111; // jalr r6, r1, 20 #r6 = 44
    	    icache[11] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 41
    	    icache[12] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 42
    	    icache[13] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 43
    	    icache[14] <= 32'b111111010101_00001_000_01000_1100111; // jalr r8, r1, -43 #r2 = 60
    	    icache[15] <= 32'b000000000100_00001_000_00111_1100111; // jalr r7, r1, 4 #r2 = 64
	    `endif
    	`ifdef TEST_BEQ
    	    icache[0] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1
    	    icache[1] <= 32'b0_000000_00001_00001_000_0100_0_1100011; // beq r1, r1, 8 # branch to 12
    	    icache[2] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r1, 1 # shouldn't happen, jumped over
    	    icache[3] <= 32'b0_000000_00001_00000_000_0100_0_1100011; // beq r0, r1, 8 # no branch
    	    icache[4] <= 32'b000000000001_00000_000_00010_0010011; // addi r2, r0, 1 #r2 = 1 
    	    icache[5] <= 32'b0_000000_00010_00001_000_0110_0_1100011; // beq r1, r2, 12 # branch to 32
    	    icache[6] <= 32'b0_000000_00010_00001_000_0110_0_1100011; // beq r1, r2, 12 # branch to 36
    	    icache[7] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r1, 1 # shouldn't happen, jumped over
    	    icache[8] <= 32'b1_111111_00001_00001_000_1100_1_1100011; // beq r1, r1, -8 # branch to 24
    	    icache[9] <= 32'b1_111111_00000_00001_000_1100_1_1100011; // beq r1, r0, -8 # no branch
    	    icache[10] <= 32'b0_000000_00010_00001_000_1010_0_1100011; // beq r1, r2, 20 # branch to 60
    	    icache[11] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1 #shouldn't happen
    	    icache[12] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1
    	    icache[13] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1
    	    icache[14] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1
    	    icache[15] <= 32'b1_111110_00010_00001_000_0010_1_1100011; // beq r1, r1, -60 #branch to 0
	    `endif
    	`ifdef TEST_BNE
    	    icache[0] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1
    	    icache[1] <= 32'b0_000000_00000_00001_001_0100_0_1100011; // bne r1, r0, 8 # branch to 12
    	    icache[2] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r1, 1 # shouldn't happen, jumped over
    	    icache[3] <= 32'b0_000000_00001_00001_001_0100_0_1100011; // bne r1, r1, 8 # no branch
    	    icache[4] <= 32'b000000000001_00000_000_00010_0010011; // addi r2, r0, 1 #r2 = 1 
    	    icache[5] <= 32'b0_000000_00000_00001_001_0110_0_1100011; // bne r1, r0, 12 # branch to 32
    	    icache[6] <= 32'b0_000000_00000_00001_001_0110_0_1100011; // bne r1, r0, 12 # branch to 36
    	    icache[7] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r1, 1 # shouldn't happen, jumped over
    	    icache[8] <= 32'b1_111111_00000_00010_001_1100_1_1100011; // bne r2, r0, -8 # branch to 24
    	    icache[9] <= 32'b1_111111_00010_00001_001_1100_1_1100011; // bne r1, r2, -8 # no branch
    	    icache[10] <= 32'b0_000000_00000_00001_001_1010_0_1100011; // bne r1, r0, 20 # branch to 60
    	    icache[11] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1 #shouldn't happen
    	    icache[12] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1
    	    icache[13] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1
    	    icache[14] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1
    	    icache[15] <= 32'b1_111110_00001_00000_001_0010_1_1100011; // bne r0, r1, -60 #branch to 0
	    `endif
    	`ifdef TEST_BLT
    	    icache[0] <= 32'b000000000010_00000_000_00001_0010011; // addi r1, r0, 2 #r1 = 2
    	    icache[1] <= 32'b000000000011_00000_000_00010_0010011; // addi r2, r0, 3 #r2 = 3
    	    icache[2] <= 32'b111111111110_00000_000_00011_0010011; // addi r3, r0, -2 #r3 = -2
    	    icache[3] <= 32'b111111111101_00000_000_00100_0010011; // addi r4, r0, -3 #r4 = -3
    	    icache[4] <= 32'b000000000001_00000_000_00000_0010011; // addi r0, r0, 1 # nop
    	    icache[5] <= 32'b0_000000_00010_00001_100_0100_0_1100011; // blt r1, r2, 8 # branch to 28
    	    icache[6] <= 32'b000000000001_00000_000_00101_0010011; // addi r5, r0, 1 # shouldn't happen, jumped over
    	    icache[7] <= 32'b0_000000_00011_00100_100_0100_0_1100011; // blt r4, r3, 8 # branch to 36
    	    icache[8] <= 32'b000000000001_00000_000_00101_0010011; // addi r5, r0, 1 # shouldn't happen, jumped over
    	    icache[9] <= 32'b0_000000_00011_00001_100_0100_0_1100011; // blt r1, r3, 8 shouldn't branch
    	    icache[10] <= 32'b0_000000_00010_00100_100_0100_0_1100011; // blt r4, r2, 8 branch to 48
    	    icache[11] <= 32'b000000000001_00000_000_00110_0010011; // addi r6, r0, 1 #r1 = 1 # r1 = 1 #shouldn't happen
    	    icache[12] <= 32'b0_000000_00000_00100_100_0100_0_1100011; // blt r4, r0, 8 branch to 56
    	    icache[13] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1
    	    icache[14] <= 32'b0_000000_00000_00010_100_0100_0_1100011; // blt r2, r0, 8 no branch
    	    icache[15] <= 32'b1_111110_00001_00100_100_0010_1_1100011; // blt r4, r1, -60 #branch to 0
	    `endif
    	`ifdef TEST_BLTU
    	    icache[0] <= 32'b000000000010_00000_000_00001_0010011; // addi r1, r0, 2 #r1 = 2
    	    icache[1] <= 32'b000000000011_00000_000_00010_0010011; // addi r2, r0, 3 #r2 = 3
    	    icache[2] <= 32'b111111111110_00000_000_00011_0010011; // addi r3, r0, -2 #r3 = -2
    	    icache[3] <= 32'b111111111101_00000_000_00100_0010011; // addi r4, r0, -3 #r4 = -3
    	    icache[4] <= 32'b000000000001_00000_000_00000_0010011; // addi r0, r0, 1 # nop
    	    icache[5] <= 32'b0_000000_00010_00001_101_0100_0_1100011; // blt r1, r2, 8 # branch to 28
    	    icache[6] <= 32'b000000000001_00000_000_00101_0010011; // addi r5, r0, 1 # shouldn't happen, jumped over
    	    icache[7] <= 32'b0_000000_00011_00100_101_0100_0_1100011; // blt r4, r3, 8 # branch to 36
    	    icache[8] <= 32'b000000000001_00000_000_00101_0010011; // addi r5, r0, 1 # shouldn't happen, jumped over
    	    icache[9] <= 32'b0_000000_00011_00001_101_0100_0_1100011; // blt r1, r3, 8 branch to 44
    	    icache[10] <= 32'b000000000001_00000_000_00110_0010011; // addi r6, r0, 1 # r1 = 1 #shouldn't happen
    	    icache[11] <= 32'b0_000000_00010_00100_101_0100_0_1100011; // blt r4, r2, 8 no branch
    	    icache[12] <= 32'b0_000000_00000_00100_101_0100_0_1100011; // blt r4, r0, 8 no branch
    	    icache[13] <= 32'b0_000000_00100_00000_101_0100_0_1100011; // blt r0, r4, 8 branch to 60
    	    icache[14] <= 32'b000000000001_00000_000_00110_0010011; // addi r6, r0, 1 # r1 = 1 #shouldn't happen
    	    icache[15] <= 32'b1_111110_00100_00001_101_0010_1_1100011; // blt r1, r4, -60 #branch to 0
	    `endif
    	`ifdef TEST_BGE
    	    icache[0] <= 32'b000000000010_00000_000_00001_0010011; // addi r1, r0, 2 #r1 = 2
    	    icache[1] <= 32'b000000000011_00000_000_00010_0010011; // addi r2, r0, 3 #r2 = 3
    	    icache[2] <= 32'b111111111110_00000_000_00011_0010011; // addi r3, r0, -2 #r3 = -2
    	    icache[3] <= 32'b111111111101_00000_000_00100_0010011; // addi r4, r0, -3 #r4 = -3
    	    icache[4] <= 32'b000000000001_00000_000_00000_0010011; // addi r0, r0, 1 # nop
    	    icache[5] <= 32'b0_000000_00001_00010_110_0100_0_1100011; // bge r2, r1, 8 # branch to 28
    	    icache[6] <= 32'b000000000001_00000_000_00101_0010011; // addi r5, r0, 1 # shouldn't happen, jumped over
    	    icache[7] <= 32'b0_000000_00100_00011_110_0100_0_1100011; // bge r3, r4, 8 # branch to 36
    	    icache[8] <= 32'b000000000001_00000_000_00101_0010011; // addi r5, r0, 1 # shouldn't happen, jumped over
    	    icache[9] <= 32'b0_000000_00001_00011_110_0100_0_1100011; // bge r3, r1, 8 shouldn't branch
    	    icache[10] <= 32'b0_000000_00100_00010_110_0100_0_1100011; // bge r2, r4, 8 branch to 48
    	    icache[11] <= 32'b000000000001_00000_000_00110_0010011; // addi r6, r0, 1 #r1 = 1 # r1 = 1 #shouldn't happen
    	    icache[12] <= 32'b0_000000_00100_00100_110_0100_0_1100011; // bge r4, r4, 8 branch to 56
    	    icache[13] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1
    	    icache[14] <= 32'b0_000000_00010_00011_110_0100_0_1100011; // bge r3, r2, 8 no branch
    	    icache[15] <= 32'b1_111110_00100_00000_110_0010_1_1100011; // bge r0, r4, -60 #branch to 0
	    `endif
    	`ifdef TEST_BGEU
    	    icache[0] <= 32'b000000000010_00000_000_00001_0010011; // addi r1, r0, 2 #r1 = 2
    	    icache[1] <= 32'b000000000011_00000_000_00010_0010011; // addi r2, r0, 3 #r2 = 3
    	    icache[2] <= 32'b111111111110_00000_000_00011_0010011; // addi r3, r0, -2 #r3 = -2
    	    icache[3] <= 32'b111111111101_00000_000_00100_0010011; // addi r4, r0, -3 #r4 = -3
    	    icache[4] <= 32'b000000000001_00000_000_00000_0010011; // addi r0, r0, 1 # nop
    	    icache[5] <= 32'b0_000000_00001_00010_111_0100_0_1100011; // bge r2, r1, 8 # branch to 28
    	    icache[6] <= 32'b000000000001_00000_000_00101_0010011; // addi r5, r0, 1 # shouldn't happen, jumped over
    	    icache[7] <= 32'b0_000000_00100_00011_111_0100_0_1100011; // bge r3, r4, 8 # branch to 36
    	    icache[8] <= 32'b000000000001_00000_000_00101_0010011; // addi r5, r0, 1 # shouldn't happen, jumped over
    	    icache[9] <= 32'b0_000000_00011_00001_111_0100_0_1100011; // bge r1, r3, 8 shouldn't branch
    	    icache[10] <= 32'b0_000000_00010_00100_111_0100_0_1100011; // bge r4, r2, 8 branch to 48
    	    icache[11] <= 32'b000000000001_00000_000_00110_0010011; // addi r6, r0, 1 #r1 = 1 # r1 = 1 #shouldn't happen
    	    icache[12] <= 32'b0_000000_00000_00100_111_0100_0_1100011; // bge r4, r0, 8 branch to 56
    	    icache[13] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 1 # r1 = 1
    	    icache[14] <= 32'b0_000000_00011_00100_111_0100_0_1100011; // bge r4, r3, 8 no branch
    	    icache[15] <= 32'b1_111110_00100_00100_111_0010_1_1100011; // bge r4, r4, -60 #branch to 0
	    `endif
    	`ifdef TEST_SW_LW_1
    	    icache[0] <= 32'b000000100000_00000_000_00001_0010011; // addi r1, r0, 32 #r1 = 32
    	    icache[1] <= 32'b000000001111_00000_000_00010_0010011; // addi r2, r0, 15 #r2 = 15
    	    icache[2] <= 32'b000011110000_00000_000_00011_0010011; // addi r3, r0, 240 #r3 = 240
    	    icache[3] <= 32'b100000000000_00000_000_00100_0010011; // addi r4, r0, -2048 #r4 = -2048
    	    icache[4] <= 32'b00000000000000001111_01010_0110111; // lui r10, 15 #r10 = 61440
    	    icache[5] <= 32'b1111111_00010_00001_010_00000_0100011; // sw r2, r1(-32) # store r2 into address 0
    	    icache[6] <= 32'b0000000_00011_00000_010_00100_0100011; // sw r3, r0(4) # store r3 into address 4
    	    icache[7] <= 32'b0000000_00100_00000_010_01000_0100011; // sw r4, r0(8) # store r4 into address 8
    	    icache[8] <= 32'b111111100000_00001_010_00101_0000011; // lw r5, r1(-32) # r5 = 15 load address 0 into r5
    	    icache[9] <= 32'b111111100100_00001_010_00110_0000011; // lw r6, r1(-28) # r6 = 240 load address 4 into r6
    	    icache[10] <= 32'b000000001000_00000_010_00111_0000011; // lw r7, r0(8) # r7 = -2048 load address 8 into r7
    	    icache[11] <= 32'b000000000100_00000_000_01000_0000011; // lb r8, r0(4) # r8 = -16 load byte at address 4 into r8
    	    icache[12] <= 32'b000000000100_00000_100_01001_0000011; // lbu r9, r0(4) # r9 = 240 load byte unsigned at address 4 into r8
    	    icache[13] <= 32'b0000000_01010_00000_010_01100_0100011; // sw r10, r0(12) # store r10 into address 12
    	    icache[14] <= 32'b000000001100_00000_001_01011_0000011; // lh r11, r0(4) # r11 = -4096 load byte at address 4 into r8
    	    icache[15] <= 32'b000000001100_00000_101_01100_0000011; // lhu r12, r0(4) # r2 = 61440 load byte at address 4 into r8
	    `endif
    	`ifdef TEST_SW_LW_2
    	    icache[0] <= 32'b111111111111_00000_000_00001_0010011; // addi r1, r0, -1 #r1 = -1
    	    icache[1] <= 32'b0000000_00001_00000_000_00000_0100011; // sb r1, r0(0) # store byte of r1 into address 0
    	    icache[2] <= 32'b0000000_00001_00000_001_00100_0100011; // sh r1, r0(4) # store half of r1 into address 4
    	    icache[3] <= 32'b000000000000_00000_000_00010_0000011; // lb r2, r0(0) # r2 = -1 load byte address 0 into r2
    	    icache[4] <= 32'b000000000100_00000_001_00011_0000011; // lh r3, r0(4) # r3 = -1 load half address 4 into r3
    	    icache[5] <= 32'b000000000000_00000_010_00100_0000011; // lw r4, r0(0) # r4 = ff load address 0 into r4
    	    icache[6] <= 32'b000000000100_00000_010_00101_0000011; // lw r5, r0(4) # r5 = ffff load address 4 into r5
    	    icache[7] <= 32'b000000000000_00000_000_00000_0010011; // nop
    	    icache[8] <= 32'b000000000000_00000_000_00000_0010011; // nop
    	    icache[9] <= 32'b000000000000_00000_000_00000_0010011; // nop
    	    icache[10] <= 32'b000000000000_00000_000_00000_0010011; // nop
    	    icache[11] <= 32'b000000000000_00000_000_00000_0010011; // nop
    	    icache[12] <= 32'b000000000000_00000_000_00000_0010011; // nop
    	    icache[13] <= 32'b000000000000_00000_000_00000_0010011; // nop
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // nop
    	    icache[15] <= 32'b000000000000_00000_000_00000_0010011; // nop
	    `endif
    	`ifdef TEST_ISSUE
    	    icache[0] <= 32'b000000000001_00000_000_00001_0010011; // addi r1, r0, 1 #r1 = 1
    	    icache[1] <= 32'b0000000_00001_00000_000_00010_1111000; // add4 v2, v0, v1 # v8-v11 = 64'h0011001100110011
    	    icache[2] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 2
    	    icache[3] <= 32'b0000000_00010_00010_000_00011_1111000; // add4 v3, v2, v2 # v12-v15 = 64'h0022002200220022
    	    icache[4] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 3
    	    icache[5] <= 32'b0000000_00010_00010_000_00011_1111001; // mult4 v3, v2, v2 # v12-v15 = 64'h0484048404840484
    	    icache[6] <= 32'b000000000001_00001_000_00001_0010011; // addi r1, r1, 1 #r1 = 4
    	    icache[7] <= 32'b0000000_00010_00010_000_00100_1111000; // add4 v4, v2, v2 # v16-v19 = 64'h0022002200220022
    	    icache[8] <= 32'b000000100000_00000_000_00010_0010011; // addi r2, r0, 32 #r2 = 32 (base address for mem)
    	    icache[9] <= 32'b000000000001_00000_000_00011_0010011; // addi r3, r0, 1 #r3 = 1 (quadword aligned stride)
    	    icache[10] <= 32'b000000000001_00010_000_00101_1111010; // load4 v5, r2(1) # v20-23 = mem[32-56]
    	    icache[11] <= 32'b000000000001_00000_000_00011_1111011; // store4 v3, r0(1) # mem[0-24] = v12-v15
    	    icache[12] <= 32'b000000000001_00010_000_00101_1111010; // load4 v5, r2(1) # v20-23 = mem[32-56]
    	    icache[13] <= 32'b000000000000_00110_000_01000_1111100; // relu4 v8, v6 # v32-35 = relu(v24-27)
    	    icache[14] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[15] <= 32'b1_111111_00000_00000_000_1110_1_1100011; // beq r0, r0, -4 # branch to 14
	    `endif
	    `ifdef TEST_MATMUL
	        // r0 is base pointer to weights1
    	    icache[0] <= 32'b00000000000000000110_00001_0110111; // lui r1, 0x00006 #r1 = 0x00006000
    	    icache[1] <= 32'b001000000000_00001_000_00001_0010011; // addi r1, r1, 0x200 #r1 = 0x00006200 //base pointer to weights2
    	    icache[2] <= 32'b00000000000000000110_00010_0110111; // lui r2, 0x00006 #r2 = 0x00006000
    	    icache[3] <= 32'b001110000000_00010_000_00010_0010011; // addi r2, r2, 0x380 #r2 = 0x00006380 //base pointer to bias1
    	    icache[4] <= 32'b00000000000000000110_00011_0110111; // lui r3, 0x00006 #r3 = 0x00006000
    	    icache[5] <= 32'b001110100000_00011_000_00011_0010011; // addi r3, r3, 0x3a0 #r3 = 0x000063a0 //base pointer to bias2
    	    icache[6] <= 32'b00000000000000001000_00100_0110111; // lui r4, 0x00008 #r4 = 0x00008000 //imagearray ptr
    	    icache[7] <= 32'b00000000000000001010_00101_0110111; // lui r5, 0x0000a #r5 = 0x0000a000 //user memory ptr
    	    icache[8] <= 32'b001100010000_00000_000_00110_0010011; // addi r6, r0, 784 #r6 = 0x310 // loop bound is 784
    	    icache[9] <= 32'b000000000000_00000_000_00111_0010011; // addi r7, r0, 0 #r7 = 0 // loop starting index is 0
    	    icache[10] <= 32'b000000000000_00100_000_01000_0010011; // addi r8, r4, 0 #r8 = 0x00008000 // r8 is now imagearray[0]
    	    icache[11] <= 32'b000011000100_01000_000_00101_1111010; // load4 v5, r8(196) # v20-23 = imagearray[0,196,392,588]
    	    icache[12] <= 32'b000000001000_01000_000_01000_0010011; // addi r8, r8, 8 #increment imagearray pointer
    	    icache[13] <= 32'b000000000000_00000_000_01001_0010011; // addi r9, r0, 0 #r9 = 0x00000000 // r9 is now weights1[0]
    	    icache[14] <= 32'b000000000100_01001_000_00110_1111010; // load4 v6, r9(4) # v24-27 = mem[0,4,8,12]
    	    icache[15] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 = 0x00000008 // r9 is now weights1[1]
    	    icache[16] <= 32'b000000000100_01001_000_00111_1111010; // load4 v7, r9(4) # v28-31 = mem[1,5,9,13]
    	    icache[17] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 = 0x00000010 // r9 is now weights1[2]
    	    icache[18] <= 32'b000000000100_01001_000_01000_1111010; // load4 v8, r9(4) # v32-35 = mem[2,6,10,14]
    	    icache[19] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 = 0x00000018 // r9 is now weights1[3]
    	    icache[20] <= 32'b000000000100_01001_000_01001_1111010; // load4 v9, r9(4) # v36-39 = mem[3,7,11,15]
    	    icache[21] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 = 0x00000020 // r9 is now weights1[4]
    	    icache[22] <= 32'b000001100000_01001_000_01001_0010011; // addi r9, r9, 96 #r9 = 0x00000080 // r9 is now weights1[16]
    	    icache[23] <= 32'b0000000_00110_00101_000_00001_1111001; // mult4 v1, v5, v6 # v4-v7 = 64'h0000000000000000
    	    icache[24] <= 32'b0000000_00111_00101_000_00010_1111001; // mult4 v2, v5, v7 # v8-v11 = 64'h0000000000000000
    	    icache[25] <= 32'b0000000_01000_00101_000_00011_1111001; // mult4 v3, v5, v8 # v12-v15 = 64'h0000000000000000
    	    icache[26] <= 32'b0000000_01001_00101_000_00100_1111001; // mult4 v4, v5, v9 # v16-v19 = 64'h0000000000000000
    	    icache[27] <= 32'b000000000100_00111_000_00111_0010011; // addi r0, r0, 0 #this should actually be r7+=4 otherwise i'm doing 1 extra loop iteration /****************loop start**********/
    	    icache[28] <= 32'b000000000100_00111_000_00111_0010011; // addi r7, r7, 4 #r7 +=4 // increment loop index
    	    icache[29] <= 32'b000011000100_01000_000_00101_1111010; // load4 v5, r8(196) # v20-23 = imagearray[1,197,393,589]
    	    icache[30] <= 32'b000000001000_01000_000_01000_0010011; // addi r8, r8, 8 #increment imagearray pointer
    	    icache[31] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[32] <= 32'b000000000100_01001_000_00110_1111010; // load4 v6, r9(4) # v24-27 = mem[0,4,8,12]
    	    icache[33] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 = 0x00000008 // r9 is now weights1[1]
    	    icache[34] <= 32'b000000000100_01001_000_00111_1111010; // load4 v7, r9(4) # v28-31 = mem[1,5,9,13]
    	    icache[35] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 = 0x00000010 // r9 is now weights1[2]
    	    icache[36] <= 32'b000000000100_01001_000_01000_1111010; // load4 v8, r9(4) # v32-35 = mem[2,6,10,14]
    	    icache[37] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 = 0x00000018 // r9 is now weights1[3]
    	    icache[38] <= 32'b000000000100_01001_000_01001_1111010; // load4 v9, r9(4) # v36-39 = mem[3,7,11,15]
    	    icache[39] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 = 0x00000020 // r9 is now weights1[4]
    	    icache[40] <= 32'b000001100000_01001_000_01001_0010011; // addi r9, r9, 96 #r9 = 0x00000080 // r9 is now weights1[16]
    	    icache[41] <= 32'b0000000_00110_00101_000_01010_1111001; // mult4 v10, v5, v6 # v40-v43 = product0
    	    icache[42] <= 32'b0000000_00111_00101_000_01011_1111001; // mult4 v11, v5, v7 # v44-v47 = product1
    	    icache[43] <= 32'b0000000_01000_00101_000_01100_1111001; // mult4 v12, v5, v8 # v48-v51 = product2
    	    icache[44] <= 32'b0000000_01001_00101_000_01101_1111001; // mult4 v13, v5, v9 # v52-v55 = product3
    	    icache[45] <= 32'b0000000_01010_00001_000_00001_1111000; // add4 v1, v1, v10 # v4-v7 accumulate
    	    icache[46] <= 32'b0000000_01011_00010_000_00010_1111000; // add4 v2, v2, v11 # v4-v7 accumulate
    	    icache[47] <= 32'b0000000_01100_00011_000_00011_1111000; // add4 v3, v3, v12 # v4-v7 accumulate
    	    icache[48] <= 32'b0000000_01101_00100_000_00100_1111000; // add4 v4, v4, v13 # v4-v7 accumulate
    	    icache[49] <= 32'b1_111101_00110_00111_100_0110_1_1100011; // blt r7, r6, 8 # branch to 32
    	    icache[50] <= 32'b000000000000_00101_000_01010_0010011; // addi r10, r5, 0 # r10 is now user memory ptr
    	    icache[51] <= 32'b000000000100_01010_000_00001_1111011; // store4 v1, r10(4) # mem[0-31] = v4=7
    	    icache[52] <= 32'b000000001000_01010_000_01010_0010011; // addi r10, r10, 8 # increment user ptr
    	    icache[53] <= 32'b000000000100_01010_000_00010_1111011; // store4 v2, r10(4) # mem[0-31] = v4=7
    	    icache[54] <= 32'b000000001000_01010_000_01010_0010011; // addi r10, r10, 8 # increment user ptr
    	    icache[55] <= 32'b000000000100_01010_000_00011_1111011; // store4 v3, r10(4) # mem[0-31] = v4=7
    	    icache[56] <= 32'b000000001000_01010_000_01010_0010011; // addi r10, r10, 8 # increment user ptr
    	    icache[57] <= 32'b000000000100_01010_000_00100_1111011; // store4 v4, r10(4) # mem[0-31] = v4=7
    	    icache[58] <= 32'b000000000001_00101_000_01110_1111010; // load4 v14, r5(1) # v56-59 = mem[0-3]
    	    icache[59] <= 32'b000000000001_00010_000_01111_1111010; // load4 v15, r2(1) # v60-63 = bias1[0-3]
    	    icache[60] <= 32'b0000000_01111_01110_000_10000_1111000; // add4 v16, v14, v15 # v64-67 bias1result
    	    icache[61] <= 32'b000000000000_10000_000_10001_1111100; // relu4 v17, v16 # v68-71 = relu(v68-71)
    	    icache[62] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop /***************first layer done****************/
    	    icache[63] <= 32'b000000100000_00101_000_01010_0010011; // addi r10, r5, 32 # r10 is now user memory ptr +32
    	    icache[64] <= 32'b000000000100_01010_000_10001_1111011; // store4 v17, r10(4) # mem[0-31] = v68-71
    	    icache[65] <= 32'b000000000001_01010_000_00100_1111010; // load4 v4, 10(1) # v16-19 = mem[32-63]
    	    icache[66] <= 32'b000000100000_00101_000_01010_0010011; // addi r10, r5, 32 # r10 is now user memory ptr +64
    	    icache[67] <= 32'b000000000000_00001_000_01001_0010011; // addi r9, r1, 0 $ r9 is weights2 ptr
    	    icache[68] <= 32'b000000000011_01001_000_00101_1111010; // load4 v5, r9(3) # v24-27 = mem[0,3,6,9]
    	    icache[69] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 += 8 // r9 is now weights2[1]
    	    icache[70] <= 32'b000000000011_01001_000_00110_1111010; // load4 v6, r9(3) # v24-27 = mem[1,4,7,10]
    	    icache[71] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 += 8 // r9 is now weights2[2]
    	    icache[72] <= 32'b000000000011_01001_000_00111_1111010; // load4 v7, r9(3) # v24-27 = mem[2,5,8,11]
    	    icache[73] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 +=8 // r9 is now weights2[3]
    	    icache[74] <= 32'b000001001000_01001_000_01001_0010011; // addi r9, r9, 72 #r9 +=72 // r9 is now weights2[3]
    	    icache[75] <= 32'b0000000_00101_00100_000_00001_1111001; // mult4 v1, v4, v5 # v4-v7 = first third
    	    icache[76] <= 32'b0000000_00110_00100_000_00010_1111001; // mult4 v2, v4, v6 # v8-v11 = second third
    	    icache[77] <= 32'b0000000_00111_00100_000_00011_1111001; // mult4 v3, v4, v7 # v12-v15 = third
    	    icache[78] <= 32'b000000010000_00000_000_00110_0010011; // addi r6, r0, 16 #r6 is outer loop index
    	    icache[79] <= 32'b000000000100_00000_000_00111_0010011; // addi r7, r0, 4 #r7 is loop counter
    	    icache[80] <= 32'b000000000001_01010_000_00100_1111010; // load4 v4, 10(1) # v16-19 = mem[32-63] //load next input matrix
    	    icache[81] <= 32'b000000100000_00101_000_01010_0010011; // addi r10, r5, 32 # r10 +=32
    	    icache[82] <= 32'b000000000011_01001_000_00101_1111010; // load4 v5, r9(3) # v24-27 = mem[0,3,6,9]
    	    icache[83] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 += 8 // r9 is now weights2[1]
    	    icache[84] <= 32'b000000000011_01001_000_00110_1111010; // load4 v6, r9(3) # v24-27 = mem[1,4,7,10]
    	    icache[85] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 += 8 // r9 is now weights2[2]
    	    icache[86] <= 32'b000000000011_01001_000_00111_1111010; // load4 v7, r9(3) # v24-27 = mem[2,5,8,11]
    	    icache[87] <= 32'b000000001000_01001_000_01001_0010011; // addi r9, r9, 8 #r9 +=8 // r9 is now weights2[3]
    	    icache[88] <= 32'b000001001000_01001_000_01001_0010011; // addi r9, r9, 72 #r9 +=72 // r9 is now weights2[3]
    	    icache[89] <= 32'b0000000_00101_00100_000_01000_1111001; // mult4 v8, v4, v5 # v32-35 = first third
    	    icache[90] <= 32'b0000000_00110_00100_000_01001_1111001; // mult4 v9, v4, v6 # v36-39 = second third
    	    icache[91] <= 32'b0000000_00111_00100_000_01010_1111001; // mult4 v10, v4, v7 # v40-43 = third
    	    icache[92] <= 32'b0000000_01000_00001_000_00001_1111000; // add4 v1, v1, v8 # accumulate first
    	    icache[93] <= 32'b0000000_01001_00010_000_00010_1111000; // add4 v2, v2, v9 # accumulate first
    	    icache[94] <= 32'b0000000_01010_00011_000_00011_1111000; // add4 v3, v3, v10 # accumulate first
    	    icache[95] <= 32'b000000000100_00111_000_00111_0010011; // addi r7, r7, 4 #r7 is loop counter
    	    icache[96] <= 32'b1_111110_00110_00111_100_0000_1_1100011; // blt r7, r6, 8 # branch to 80
    	    icache[97] <= 32'b000000000000_00101_000_01010_0010011; // addi r10, r5, 0 # r10 is now user memory ptr
    	    icache[98] <= 32'b000000100000_01010_000_01010_0010011; // addi r10, r10, 32 # increment user ptr by 32 (next 32 byte segment)
    	    icache[99] <= 32'b000000000100_01010_000_00001_1111011; // store4 v1, r10(4) # mem[0-31] = v4=7
    	    icache[100] <= 32'b000000001000_01010_000_01010_0010011; // addi r10, r10, 8 # increment user ptr by 8
    	    icache[101] <= 32'b000000000100_01010_000_00010_1111011; // store4 v2, r10(4) # mem[0-31] = v4=7
    	    icache[102] <= 32'b000000001000_01010_000_01010_0010011; // addi r10, r10, 8 # increment user ptr by 8
    	    icache[103] <= 32'b000000000100_01010_000_00011_1111011; // store4 v3, r10(4) # mem[0-31] = v4=7
    	    icache[104] <= 32'b000000100000_00101_000_01010_0010011; // addi r10, r5, 32 # r10 is now user memory ptr at second 32bytes
    	    icache[105] <= 32'b000000000001_01010_000_01011_1111010; // load4 v11, r5(1) # v44-47 = mem[4-7]
    	    icache[106] <= 32'b000000000001_00011_000_01100_1111010; // load4 v12, r3(1) # v48-51 = bias2[0-3]
    	    icache[107] <= 32'b0000000_01100_01011_000_01101_1111000; // add4 v13, v11, v12 # v52-55 finalresult
    	    icache[108] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[109] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[110] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[111] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[112] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[113] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[114] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[115] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[116] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[117] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[118] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[119] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[120] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[121] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[122] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[123] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[124] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[125] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[126] <= 32'b000000000000_00000_000_00000_0010011; // addi r0, r0, 0 #nop
    	    icache[127] <= 32'b1_111111_00000_00000_000_1110_1_1100011; // beq r0, r0, -4 # branch to 126
	    `endif
    	end else begin
    	// do nothing
    	end
    end

endmodule
