module dcache_image(address, read, data_out, valid, CLK, RST);
    parameter WIDTH = 32;
    parameter VEC_WIDTH = 64;
    reg [VEC_WIDTH-1:0] dcache [1023:0];
    
    input wire [WIDTH-1:0] address;
    input wire read;
    output wire [VEC_WIDTH-1:0] data_out;
    output wire valid;
    input CLK, RST;
    
    assign valid = 1'b1;
    
    wire [9:0] index = address[12:3];
    
    //always do this no matter what (read always active basically)
    assign data_out = dcache[index];
    
    initial begin
        dcache[0] <= 64'h0000000000000000;
        dcache[1] <= 64'h0000000000000000;
        dcache[2] <= 64'h0000000000000000;
        dcache[3] <= 64'h0000000000000000;
        dcache[4] <= 64'h0000000000000000;
        dcache[5] <= 64'h0000000000000000;
        dcache[6] <= 64'h0000000000000000;
        dcache[7] <= 64'h0000000000000000;
        dcache[8] <= 64'h0000000000000000;
        dcache[9] <= 64'h0000000000000000;
        dcache[10] <= 64'h0000000000000000;
        dcache[11] <= 64'h0000000000000000;
        dcache[12] <= 64'h0000000000000000;
        dcache[13] <= 64'h0000000000000000;
        dcache[14] <= 64'h0000000000000000;
        dcache[15] <= 64'h0000000000000000;
        dcache[16] <= 64'h0000000000000000;
        dcache[17] <= 64'h0000000000000000;
        dcache[18] <= 64'h0000000000000000;
        dcache[19] <= 64'h0000000000000000;
        dcache[20] <= 64'h0000000000000000;
        dcache[21] <= 64'h0000000000000000;
        dcache[22] <= 64'h0000000000000000;
        dcache[23] <= 64'h0000000000000000;
        dcache[24] <= 64'h0000000000000000;
        dcache[25] <= 64'h0000000000000000;
        dcache[26] <= 64'h0000000000000000;
        dcache[27] <= 64'h0000000000000000;
        dcache[28] <= 64'h0000000000000000;
        dcache[29] <= 64'h0000000000000000;
        dcache[30] <= 64'h0000000000000000;
        dcache[31] <= 64'h0000000000000000;
        dcache[32] <= 64'h0000000000000000;
        dcache[33] <= 64'h0000000000000000;
        dcache[34] <= 64'h0000000000000000;
        dcache[35] <= 64'h0000000000000000;
        dcache[36] <= 64'h0000000000000000;
        dcache[37] <= 64'h0000000000c80383;
        dcache[38] <= 64'h0000000000000000;
        dcache[39] <= 64'h0000000000000119;
        dcache[40] <= 64'h0074000000000000;
        dcache[41] <= 64'h0000000000000000;
        dcache[42] <= 64'h0000000000000000;
        dcache[43] <= 64'h0000000000000000;
        dcache[44] <= 64'h0000000001e5039f;
        dcache[45] <= 64'h0000000000000000;
        dcache[46] <= 64'h0000000000000252;
        dcache[47] <= 64'h02a2000000000000;
        dcache[48] <= 64'h0000000000000000;
        dcache[49] <= 64'h0000000000000000;
        dcache[50] <= 64'h0000000000000000;
        dcache[51] <= 64'h00000010030f039f;
        dcache[52] <= 64'h0000000000000000;
        dcache[53] <= 64'h0000000000000181;
        dcache[54] <= 64'h034b002c00000000;
        dcache[55] <= 64'h0000000000000000;
        dcache[56] <= 64'h0000000000000000;
        dcache[57] <= 64'h0000000000000000;
        dcache[58] <= 64'h0000011503f3021a;
        dcache[59] <= 64'h0000000000000000;
        dcache[60] <= 64'h00000000000001c9;
        dcache[61] <= 64'h03f3005400000000;
        dcache[62] <= 64'h0000000000000000;
        dcache[63] <= 64'h0000000000000000;
        dcache[64] <= 64'h0000000000000000;
        dcache[65] <= 64'h00b403b303670030;
        dcache[66] <= 64'h0000000000000000;
        dcache[67] <= 64'h0000000000000303;
        dcache[68] <= 64'h03f3005400000000;
        dcache[69] <= 64'h0000000000000000;
        dcache[70] <= 64'h0000000000000000;
        dcache[71] <= 64'h0000000000000000;
        dcache[72] <= 64'h02a203df00d40000;
        dcache[73] <= 64'h0000000000000000;
        dcache[74] <= 64'h0000000000480400;
        dcache[75] <= 64'h03f7005400000000;
        dcache[76] <= 64'h0000000000000000;
        dcache[77] <= 64'h0000000000000000;
        dcache[78] <= 64'h0000000000000151;
        dcache[79] <= 64'h03cb034f00000000;
        dcache[80] <= 64'h0000000000000000;
        dcache[81] <= 64'h00000000023603f7;
        dcache[82] <= 64'h02f6001400000000;
        dcache[83] <= 64'h0000000000000000;
        dcache[84] <= 64'h0000000000000000;
        dcache[85] <= 64'h00000000000002a6;
        dcache[86] <= 64'h03f301a900000000;
        dcache[87] <= 64'h0000000000000000;
        dcache[88] <= 64'h0000008003a303eb;
        dcache[89] <= 64'h0109000000000000;
        dcache[90] <= 64'h0000000000000000;
        dcache[91] <= 64'h0000000000000000;
        dcache[92] <= 64'h00000000003c0387;
        dcache[93] <= 64'h03f3000000000000;
        dcache[94] <= 64'h0000000000000000;
        dcache[95] <= 64'h0000021a03f3034f;
        dcache[96] <= 64'h0000000000000000;
        dcache[97] <= 64'h0000000000000000;
        dcache[98] <= 64'h0000000000000000;
        dcache[99] <= 64'h00000000005803f3;
        dcache[100] <= 64'h0292000000000000;
        dcache[101] <= 64'h0000000000000000;
        dcache[102] <= 64'h000002a603f3029e;
        dcache[103] <= 64'h0000000000000000;
        dcache[104] <= 64'h0000000000000000;
        dcache[105] <= 64'h0000000000000000;
        dcache[106] <= 64'h0000000000240333;
        dcache[107] <= 64'h0347004800000000;
        dcache[108] <= 64'h0000000000000000;
        dcache[109] <= 64'h005803f703f701ad;
        dcache[110] <= 64'h0000000000000000;
        dcache[111] <= 64'h0000000000000000;
        dcache[112] <= 64'h0000000000000000;
        dcache[113] <= 64'h00000000000002a6;
        dcache[114] <= 64'h03f3031f01550155;
        dcache[115] <= 64'h0155015502060292;
        dcache[116] <= 64'h030f03f303f301a9;
        dcache[117] <= 64'h0000000000000000;
        dcache[118] <= 64'h0000000000000000;
        dcache[119] <= 64'h0000000000000000;
        dcache[120] <= 64'h00000000000000a4;
        dcache[121] <= 64'h02aa03d703f303f3;
        dcache[122] <= 64'h03f303f303a3039f;
        dcache[123] <= 64'h03ef03f303f30024;
        dcache[124] <= 64'h0000000000000000;
        dcache[125] <= 64'h0000000000000000;
        dcache[126] <= 64'h0000000000000000;
        dcache[127] <= 64'h0000000000000000;
        dcache[128] <= 64'h000000c401510151;
        dcache[129] <= 64'h0151015100000000;
        dcache[130] <= 64'h028603f303f30000;
        dcache[131] <= 64'h0000000000000000;
        dcache[132] <= 64'h0000000000000000;
        dcache[133] <= 64'h0000000000000000;
        dcache[134] <= 64'h0000000000000000;
        dcache[135] <= 64'h0000000000000000;
        dcache[136] <= 64'h0000000000000000;
        dcache[137] <= 64'h01fd03f303f300b4;
        dcache[138] <= 64'h0000000000000000;
        dcache[139] <= 64'h0000000000000000;
        dcache[140] <= 64'h0000000000000000;
        dcache[141] <= 64'h0000000000000000;
        dcache[142] <= 64'h0000000000000000;
        dcache[143] <= 64'h0000000000000000;
        dcache[144] <= 64'h020203f703f70000;
        dcache[145] <= 64'h0000000000000000;
        dcache[146] <= 64'h0000000000000000;
        dcache[147] <= 64'h0000000000000000;
        dcache[148] <= 64'h0000000000000000;
        dcache[149] <= 64'h0000000000000000;
        dcache[150] <= 64'h0000000000000000;
        dcache[151] <= 64'h01fd03f303f30000;
        dcache[152] <= 64'h0000000000000000;
        dcache[153] <= 64'h0000000000000000;
        dcache[154] <= 64'h0000000000000000;
        dcache[155] <= 64'h0000000000000000;
        dcache[156] <= 64'h0000000000000000;
        dcache[157] <= 64'h0000000000000000;
        dcache[158] <= 64'h021e03f303d30000;
        dcache[159] <= 64'h0000000000000000;
        dcache[160] <= 64'h0000000000000000;
        dcache[161] <= 64'h0000000000000000;
        dcache[162] <= 64'h0000000000000000;
        dcache[163] <= 64'h0000000000000000;
        dcache[164] <= 64'h0000000000000000;
        dcache[165] <= 64'h03a303b301bd0000;
        dcache[166] <= 64'h0000000000000000;
        dcache[167] <= 64'h0000000000000000;
        dcache[168] <= 64'h0000000000000000;
        dcache[169] <= 64'h0000000000000000;
        dcache[170] <= 64'h0000000000000000;
        dcache[171] <= 64'h0000000000000000;
        dcache[172] <= 64'h02ce010900000000;
        dcache[173] <= 64'h0000000000000000;
        dcache[174] <= 64'h0000000000000000;
        dcache[175] <= 64'h0000000000000000;
        dcache[176] <= 64'h0000000000000000;
        dcache[177] <= 64'h0000000000000000;
        dcache[178] <= 64'h0000000000000000;
        dcache[179] <= 64'h0000000000000000;
        dcache[180] <= 64'h0000000000000000;
        dcache[181] <= 64'h0000000000000000;
        dcache[182] <= 64'h0000000000000000;
        dcache[183] <= 64'h0000000000000000;
        dcache[184] <= 64'h0000000000000000;
        dcache[185] <= 64'h0000000000000000;
        dcache[186] <= 64'h0000000000000000;
        dcache[187] <= 64'h0000000000000000;
        dcache[188] <= 64'h0000000000000000;
        dcache[189] <= 64'h0000000000000000;
        dcache[190] <= 64'h0000000000000000;
        dcache[191] <= 64'h0000000000000000;
        dcache[192] <= 64'h0000000000000000;
        dcache[193] <= 64'h0000000000000000;
        dcache[194] <= 64'h0000000000000000;
        dcache[195] <= 64'h0000000000000000;
        dcache[196] <= 64'h0000000000000000;
        dcache[197] <= 64'h0000000000000000;
        dcache[198] <= 64'h0000000000000000;
        dcache[199] <= 64'h0000000000000000;
        dcache[200] <= 64'h0000000000000000;
        dcache[201] <= 64'h0000000000000000;
        dcache[202] <= 64'h0000000000000000;
        dcache[203] <= 64'h0000000000000000;
        dcache[204] <= 64'h0000000000000000;
        dcache[205] <= 64'h0000000000000000;
        dcache[206] <= 64'h0000000000000000;
        dcache[207] <= 64'h0000000000000000;
        dcache[208] <= 64'h0000000000000000;
        dcache[209] <= 64'h0000000000000000;
        dcache[210] <= 64'h0000000000000000;
        dcache[211] <= 64'h0000000000000000;
        dcache[212] <= 64'h0000000000000000;
        dcache[213] <= 64'h0000000000000000;
        dcache[214] <= 64'h0000000000000000;
        dcache[215] <= 64'h0000000000000000;
        dcache[216] <= 64'h0000000000000000;
        dcache[217] <= 64'h0000000000000000;
        dcache[218] <= 64'h0000000000000000;
        dcache[219] <= 64'h0000000000000000;
        dcache[220] <= 64'h0000000000000000;
        dcache[221] <= 64'h0000000000000000;
        dcache[222] <= 64'h0000000000000000;
        dcache[223] <= 64'h0000000000000000;
        dcache[224] <= 64'h0000000000000000;
        dcache[225] <= 64'h0000000000000000;
        dcache[226] <= 64'h0000000000000000;
        dcache[227] <= 64'h0000000000000000;
        dcache[228] <= 64'h0000000000000000;
        dcache[229] <= 64'h0000000000000000;
        dcache[230] <= 64'h0000000000000000;
        dcache[231] <= 64'h0000000000000000;
        dcache[232] <= 64'h0000000000000000;
        dcache[233] <= 64'h0000000000000000;
        dcache[234] <= 64'h0000000000000000;
        dcache[235] <= 64'h0000000000000000;
        dcache[236] <= 64'h0000000000000000;
        dcache[237] <= 64'h0000000000000000;
        dcache[238] <= 64'h0000000000000000;
        dcache[239] <= 64'h0000000000000000;
        dcache[240] <= 64'h0000000000000000;
        dcache[241] <= 64'h0000000000000000;
        dcache[242] <= 64'h0000000000000000;
        dcache[243] <= 64'h0000000000000000;
        dcache[244] <= 64'h0000000000000000;
        dcache[245] <= 64'h0000000000000000;
        dcache[246] <= 64'h0000000000000000;
        dcache[247] <= 64'h0000000000000000;
        dcache[248] <= 64'h0000000000000000;
        dcache[249] <= 64'h0000000000000000;
        dcache[250] <= 64'h0000000000000000;
        dcache[251] <= 64'h0000000000000000;
        dcache[252] <= 64'h0000000000000000;
        dcache[253] <= 64'h0000000000000000;
        dcache[254] <= 64'h0000000000000000;
        dcache[255] <= 64'h0000000000000000;
        dcache[256] <= 64'h0000000000000000;
        dcache[257] <= 64'h0000000000000000;
        dcache[258] <= 64'h0000000000000000;
        dcache[259] <= 64'h0000000000000000;
        dcache[260] <= 64'h0000000000000000;
        dcache[261] <= 64'h0000000000000000;
        dcache[262] <= 64'h0000000000000000;
        dcache[263] <= 64'h0000000000000000;
        dcache[264] <= 64'h0000000000000000;
        dcache[265] <= 64'h0000000000000000;
        dcache[266] <= 64'h0000000000000000;
        dcache[267] <= 64'h0000000000000000;
        dcache[268] <= 64'h0000000000000000;
        dcache[269] <= 64'h0000000000000000;
        dcache[270] <= 64'h0000000000000000;
        dcache[271] <= 64'h0000000000000000;
        dcache[272] <= 64'h0000000000000000;
        dcache[273] <= 64'h0000000000000000;
        dcache[274] <= 64'h0000000000000000;
        dcache[275] <= 64'h0000000000000000;
        dcache[276] <= 64'h0000000000000000;
        dcache[277] <= 64'h0000000000000000;
        dcache[278] <= 64'h0000000000000000;
        dcache[279] <= 64'h0000000000000000;
        dcache[280] <= 64'h0000000000000000;
        dcache[281] <= 64'h0000000000000000;
        dcache[282] <= 64'h0000000000000000;
        dcache[283] <= 64'h0000000000000000;
        dcache[284] <= 64'h0000000000000000;
        dcache[285] <= 64'h0000000000000000;
        dcache[286] <= 64'h0000000000000000;
        dcache[287] <= 64'h0000000000000000;
        dcache[288] <= 64'h0000000000000000;
        dcache[289] <= 64'h0000000000000000;
        dcache[290] <= 64'h0000000000000000;
        dcache[291] <= 64'h0000000000000000;
        dcache[292] <= 64'h0000000000000000;
        dcache[293] <= 64'h0000000000000000;
        dcache[294] <= 64'h0000000000000000;
        dcache[295] <= 64'h0000000000000000;
        dcache[296] <= 64'h0000000000000000;
        dcache[297] <= 64'h0000000000000000;
        dcache[298] <= 64'h0000000000000000;
        dcache[299] <= 64'h0000000000000000;
        dcache[300] <= 64'h0000000000000000;
        dcache[301] <= 64'h0000000000000000;
        dcache[302] <= 64'h0000000000000000;
        dcache[303] <= 64'h0000000000000000;
        dcache[304] <= 64'h0000000000000000;
        dcache[305] <= 64'h0000000000000000;
        dcache[306] <= 64'h0000000000000000;
        dcache[307] <= 64'h0000000000000000;
        dcache[308] <= 64'h0000000000000000;
        dcache[309] <= 64'h0000000000000000;
        dcache[310] <= 64'h0000000000000000;
        dcache[311] <= 64'h0000000000000000;
        dcache[312] <= 64'h0000000000000000;
        dcache[313] <= 64'h0000000000000000;
        dcache[314] <= 64'h0000000000000000;
        dcache[315] <= 64'h0000000000000000;
        dcache[316] <= 64'h0000000000000000;
        dcache[317] <= 64'h0000000000000000;
        dcache[318] <= 64'h0000000000000000;
        dcache[319] <= 64'h0000000000000000;
        dcache[320] <= 64'h0000000000000000;
        dcache[321] <= 64'h0000000000000000;
        dcache[322] <= 64'h0000000000000000;
        dcache[323] <= 64'h0000000000000000;
        dcache[324] <= 64'h0000000000000000;
        dcache[325] <= 64'h0000000000000000;
        dcache[326] <= 64'h0000000000000000;
        dcache[327] <= 64'h0000000000000000;
        dcache[328] <= 64'h0000000000000000;
        dcache[329] <= 64'h0000000000000000;
        dcache[330] <= 64'h0000000000000000;
        dcache[331] <= 64'h0000000000000000;
        dcache[332] <= 64'h0000000000000000;
        dcache[333] <= 64'h0000000000000000;
        dcache[334] <= 64'h0000000000000000;
        dcache[335] <= 64'h0000000000000000;
        dcache[336] <= 64'h0000000000000000;
        dcache[337] <= 64'h0000000000000000;
        dcache[338] <= 64'h0000000000000000;
        dcache[339] <= 64'h0000000000000000;
        dcache[340] <= 64'h0000000000000000;
        dcache[341] <= 64'h0000000000000000;
        dcache[342] <= 64'h0000000000000000;
        dcache[343] <= 64'h0000000000000000;
        dcache[344] <= 64'h0000000000000000;
        dcache[345] <= 64'h0000000000000000;
        dcache[346] <= 64'h0000000000000000;
        dcache[347] <= 64'h0000000000000000;
        dcache[348] <= 64'h0000000000000000;
        dcache[349] <= 64'h0000000000000000;
        dcache[350] <= 64'h0000000000000000;
        dcache[351] <= 64'h0000000000000000;
        dcache[352] <= 64'h0000000000000000;
        dcache[353] <= 64'h0000000000000000;
        dcache[354] <= 64'h0000000000000000;
        dcache[355] <= 64'h0000000000000000;
        dcache[356] <= 64'h0000000000000000;
        dcache[357] <= 64'h0000000000000000;
        dcache[358] <= 64'h0000000000000000;
        dcache[359] <= 64'h0000000000000000;
        dcache[360] <= 64'h0000000000000000;
        dcache[361] <= 64'h0000000000000000;
        dcache[362] <= 64'h0000000000000000;
        dcache[363] <= 64'h0000000000000000;
        dcache[364] <= 64'h0000000000000000;
        dcache[365] <= 64'h0000000000000000;
        dcache[366] <= 64'h0000000000000000;
        dcache[367] <= 64'h0000000000000000;
        dcache[368] <= 64'h0000000000000000;
        dcache[369] <= 64'h0000000000000000;
        dcache[370] <= 64'h0000000000000000;
        dcache[371] <= 64'h0000000000000000;
        dcache[372] <= 64'h0000000000000000;
        dcache[373] <= 64'h0000000000000000;
        dcache[374] <= 64'h0000000000000000;
        dcache[375] <= 64'h0000000000000000;
        dcache[376] <= 64'h0000000000000000;
        dcache[377] <= 64'h0000000000000000;
        dcache[378] <= 64'h0000000000000000;
        dcache[379] <= 64'h0000000000000000;
        dcache[380] <= 64'h0000000000000000;
        dcache[381] <= 64'h0000000000000000;
        dcache[382] <= 64'h0000000000000000;
        dcache[383] <= 64'h0000000000000000;
        dcache[384] <= 64'h0000000000000000;
        dcache[385] <= 64'h0000000000000000;
        dcache[386] <= 64'h0000000000000000;
        dcache[387] <= 64'h0000000000000000;
        dcache[388] <= 64'h0000000000000000;
        dcache[389] <= 64'h0000000000000000;
        dcache[390] <= 64'h0000000000000000;
        dcache[391] <= 64'h0000000000000000;
        dcache[392] <= 64'h0000000000000000;
        dcache[393] <= 64'h0000000000000000;
        dcache[394] <= 64'h0000000000000000;
        dcache[395] <= 64'h0000000000000000;
        dcache[396] <= 64'h0000000000000000;
        dcache[397] <= 64'h0000000000000000;
        dcache[398] <= 64'h0000000000000000;
        dcache[399] <= 64'h0000000000000000;
        dcache[400] <= 64'h0000000000000000;
        dcache[401] <= 64'h0000000000000000;
        dcache[402] <= 64'h0000000000000000;
        dcache[403] <= 64'h0000000000000000;
        dcache[404] <= 64'h0000000000000000;
        dcache[405] <= 64'h0000000000000000;
        dcache[406] <= 64'h0000000000000000;
        dcache[407] <= 64'h0000000000000000;
        dcache[408] <= 64'h0000000000000000;
        dcache[409] <= 64'h0000000000000000;
        dcache[410] <= 64'h0000000000000000;
        dcache[411] <= 64'h0000000000000000;
        dcache[412] <= 64'h0000000000000000;
        dcache[413] <= 64'h0000000000000000;
        dcache[414] <= 64'h0000000000000000;
        dcache[415] <= 64'h0000000000000000;
        dcache[416] <= 64'h0000000000000000;
        dcache[417] <= 64'h0000000000000000;
        dcache[418] <= 64'h0000000000000000;
        dcache[419] <= 64'h0000000000000000;
        dcache[420] <= 64'h0000000000000000;
        dcache[421] <= 64'h0000000000000000;
        dcache[422] <= 64'h0000000000000000;
        dcache[423] <= 64'h0000000000000000;
        dcache[424] <= 64'h0000000000000000;
        dcache[425] <= 64'h0000000000000000;
        dcache[426] <= 64'h0000000000000000;
        dcache[427] <= 64'h0000000000000000;
        dcache[428] <= 64'h0000000000000000;
        dcache[429] <= 64'h0000000000000000;
        dcache[430] <= 64'h0000000000000000;
        dcache[431] <= 64'h0000000000000000;
        dcache[432] <= 64'h0000000000000000;
        dcache[433] <= 64'h0000000000000000;
        dcache[434] <= 64'h0000000000000000;
        dcache[435] <= 64'h0000000000000000;
        dcache[436] <= 64'h0000000000000000;
        dcache[437] <= 64'h0000000000000000;
        dcache[438] <= 64'h0000000000000000;
        dcache[439] <= 64'h0000000000000000;
        dcache[440] <= 64'h0000000000000000;
        dcache[441] <= 64'h0000000000000000;
        dcache[442] <= 64'h0000000000000000;
        dcache[443] <= 64'h0000000000000000;
        dcache[444] <= 64'h0000000000000000;
        dcache[445] <= 64'h0000000000000000;
        dcache[446] <= 64'h0000000000000000;
        dcache[447] <= 64'h0000000000000000;
        dcache[448] <= 64'h0000000000000000;
        dcache[449] <= 64'h0000000000000000;
        dcache[450] <= 64'h0000000000000000;
        dcache[451] <= 64'h0000000000000000;
        dcache[452] <= 64'h0000000000000000;
        dcache[453] <= 64'h0000000000000000;
        dcache[454] <= 64'h0000000000000000;
        dcache[455] <= 64'h0000000000000000;
        dcache[456] <= 64'h0000000000000000;
        dcache[457] <= 64'h0000000000000000;
        dcache[458] <= 64'h0000000000000000;
        dcache[459] <= 64'h0000000000000000;
        dcache[460] <= 64'h0000000000000000;
        dcache[461] <= 64'h0000000000000000;
        dcache[462] <= 64'h0000000000000000;
        dcache[463] <= 64'h0000000000000000;
        dcache[464] <= 64'h0000000000000000;
        dcache[465] <= 64'h0000000000000000;
        dcache[466] <= 64'h0000000000000000;
        dcache[467] <= 64'h0000000000000000;
        dcache[468] <= 64'h0000000000000000;
        dcache[469] <= 64'h0000000000000000;
        dcache[470] <= 64'h0000000000000000;
        dcache[471] <= 64'h0000000000000000;
        dcache[472] <= 64'h0000000000000000;
        dcache[473] <= 64'h0000000000000000;
        dcache[474] <= 64'h0000000000000000;
        dcache[475] <= 64'h0000000000000000;
        dcache[476] <= 64'h0000000000000000;
        dcache[477] <= 64'h0000000000000000;
        dcache[478] <= 64'h0000000000000000;
        dcache[479] <= 64'h0000000000000000;
        dcache[480] <= 64'h0000000000000000;
        dcache[481] <= 64'h0000000000000000;
        dcache[482] <= 64'h0000000000000000;
        dcache[483] <= 64'h0000000000000000;
        dcache[484] <= 64'h0000000000000000;
        dcache[485] <= 64'h0000000000000000;
        dcache[486] <= 64'h0000000000000000;
        dcache[487] <= 64'h0000000000000000;
        dcache[488] <= 64'h0000000000000000;
        dcache[489] <= 64'h0000000000000000;
        dcache[490] <= 64'h0000000000000000;
        dcache[491] <= 64'h0000000000000000;
        dcache[492] <= 64'h0000000000000000;
        dcache[493] <= 64'h0000000000000000;
        dcache[494] <= 64'h0000000000000000;
        dcache[495] <= 64'h0000000000000000;
        dcache[496] <= 64'h0000000000000000;
        dcache[497] <= 64'h0000000000000000;
        dcache[498] <= 64'h0000000000000000;
        dcache[499] <= 64'h0000000000000000;
        dcache[500] <= 64'h0000000000000000;
        dcache[501] <= 64'h0000000000000000;
        dcache[502] <= 64'h0000000000000000;
        dcache[503] <= 64'h0000000000000000;
        dcache[504] <= 64'h0000000000000000;
        dcache[505] <= 64'h0000000000000000;
        dcache[506] <= 64'h0000000000000000;
        dcache[507] <= 64'h0000000000000000;
        dcache[508] <= 64'h0000000000000000;
        dcache[509] <= 64'h0000000000000000;
        dcache[510] <= 64'h0000000000000000;
        dcache[511] <= 64'h0000000000000000;
        dcache[512] <= 64'h0000000000000000;
        dcache[513] <= 64'h0000000000000000;
        dcache[514] <= 64'h0000000000000000;
        dcache[515] <= 64'h0000000000000000;
        dcache[516] <= 64'h0000000000000000;
        dcache[517] <= 64'h0000000000000000;
        dcache[518] <= 64'h0000000000000000;
        dcache[519] <= 64'h0000000000000000;
        dcache[520] <= 64'h0000000000000000;
        dcache[521] <= 64'h0000000000000000;
        dcache[522] <= 64'h0000000000000000;
        dcache[523] <= 64'h0000000000000000;
        dcache[524] <= 64'h0000000000000000;
        dcache[525] <= 64'h0000000000000000;
        dcache[526] <= 64'h0000000000000000;
        dcache[527] <= 64'h0000000000000000;
        dcache[528] <= 64'h0000000000000000;
        dcache[529] <= 64'h0000000000000000;
        dcache[530] <= 64'h0000000000000000;
        dcache[531] <= 64'h0000000000000000;
        dcache[532] <= 64'h0000000000000000;
        dcache[533] <= 64'h0000000000000000;
        dcache[534] <= 64'h0000000000000000;
        dcache[535] <= 64'h0000000000000000;
        dcache[536] <= 64'h0000000000000000;
        dcache[537] <= 64'h0000000000000000;
        dcache[538] <= 64'h0000000000000000;
        dcache[539] <= 64'h0000000000000000;
        dcache[540] <= 64'h0000000000000000;
        dcache[541] <= 64'h0000000000000000;
        dcache[542] <= 64'h0000000000000000;
        dcache[543] <= 64'h0000000000000000;
        dcache[544] <= 64'h0000000000000000;
        dcache[545] <= 64'h0000000000000000;
        dcache[546] <= 64'h0000000000000000;
        dcache[547] <= 64'h0000000000000000;
        dcache[548] <= 64'h0000000000000000;
        dcache[549] <= 64'h0000000000000000;
        dcache[550] <= 64'h0000000000000000;
        dcache[551] <= 64'h0000000000000000;
        dcache[552] <= 64'h0000000000000000;
        dcache[553] <= 64'h0000000000000000;
        dcache[554] <= 64'h0000000000000000;
        dcache[555] <= 64'h0000000000000000;
        dcache[556] <= 64'h0000000000000000;
        dcache[557] <= 64'h0000000000000000;
        dcache[558] <= 64'h0000000000000000;
        dcache[559] <= 64'h0000000000000000;
        dcache[560] <= 64'h0000000000000000;
        dcache[561] <= 64'h0000000000000000;
        dcache[562] <= 64'h0000000000000000;
        dcache[563] <= 64'h0000000000000000;
        dcache[564] <= 64'h0000000000000000;
        dcache[565] <= 64'h0000000000000000;
        dcache[566] <= 64'h0000000000000000;
        dcache[567] <= 64'h0000000000000000;
        dcache[568] <= 64'h0000000000000000;
        dcache[569] <= 64'h0000000000000000;
        dcache[570] <= 64'h0000000000000000;
        dcache[571] <= 64'h0000000000000000;
        dcache[572] <= 64'h0000000000000000;
        dcache[573] <= 64'h0000000000000000;
        dcache[574] <= 64'h0000000000000000;
        dcache[575] <= 64'h0000000000000000;
        dcache[576] <= 64'h0000000000000000;
        dcache[577] <= 64'h0000000000000000;
        dcache[578] <= 64'h0000000000000000;
        dcache[579] <= 64'h0000000000000000;
        dcache[580] <= 64'h0000000000000000;
        dcache[581] <= 64'h0000000000000000;
        dcache[582] <= 64'h0000000000000000;
        dcache[583] <= 64'h0000000000000000;
        dcache[584] <= 64'h0000000000000000;
        dcache[585] <= 64'h0000000000000000;
        dcache[586] <= 64'h0000000000000000;
        dcache[587] <= 64'h0000000000000000;
        dcache[588] <= 64'h0000000000000000;
        dcache[589] <= 64'h0000000000000000;
        dcache[590] <= 64'h0000000000000000;
        dcache[591] <= 64'h0000000000000000;
        dcache[592] <= 64'h0000000000000000;
        dcache[593] <= 64'h0000000000000000;
        dcache[594] <= 64'h0000000000000000;
        dcache[595] <= 64'h0000000000000000;
        dcache[596] <= 64'h0000000000000000;
        dcache[597] <= 64'h0000000000000000;
        dcache[598] <= 64'h0000000000000000;
        dcache[599] <= 64'h0000000000000000;
        dcache[600] <= 64'h0000000000000000;
        dcache[601] <= 64'h0000000000000000;
        dcache[602] <= 64'h0000000000000000;
        dcache[603] <= 64'h0000000000000000;
        dcache[604] <= 64'h0000000000000000;
        dcache[605] <= 64'h0000000000000000;
        dcache[606] <= 64'h0000000000000000;
        dcache[607] <= 64'h0000000000000000;
        dcache[608] <= 64'h0000000000000000;
        dcache[609] <= 64'h0000000000000000;
        dcache[610] <= 64'h0000000000000000;
        dcache[611] <= 64'h0000000000000000;
        dcache[612] <= 64'h0000000000000000;
        dcache[613] <= 64'h0000000000000000;
        dcache[614] <= 64'h0000000000000000;
        dcache[615] <= 64'h0000000000000000;
        dcache[616] <= 64'h0000000000000000;
        dcache[617] <= 64'h0000000000000000;
        dcache[618] <= 64'h0000000000000000;
        dcache[619] <= 64'h0000000000000000;
        dcache[620] <= 64'h0000000000000000;
        dcache[621] <= 64'h0000000000000000;
        dcache[622] <= 64'h0000000000000000;
        dcache[623] <= 64'h0000000000000000;
        dcache[624] <= 64'h0000000000000000;
        dcache[625] <= 64'h0000000000000000;
        dcache[626] <= 64'h0000000000000000;
        dcache[627] <= 64'h0000000000000000;
        dcache[628] <= 64'h0000000000000000;
        dcache[629] <= 64'h0000000000000000;
        dcache[630] <= 64'h0000000000000000;
        dcache[631] <= 64'h0000000000000000;
        dcache[632] <= 64'h0000000000000000;
        dcache[633] <= 64'h0000000000000000;
        dcache[634] <= 64'h0000000000000000;
        dcache[635] <= 64'h0000000000000000;
        dcache[636] <= 64'h0000000000000000;
        dcache[637] <= 64'h0000000000000000;
        dcache[638] <= 64'h0000000000000000;
        dcache[639] <= 64'h0000000000000000;
        dcache[640] <= 64'h0000000000000000;
        dcache[641] <= 64'h0000000000000000;
        dcache[642] <= 64'h0000000000000000;
        dcache[643] <= 64'h0000000000000000;
        dcache[644] <= 64'h0000000000000000;
        dcache[645] <= 64'h0000000000000000;
        dcache[646] <= 64'h0000000000000000;
        dcache[647] <= 64'h0000000000000000;
        dcache[648] <= 64'h0000000000000000;
        dcache[649] <= 64'h0000000000000000;
        dcache[650] <= 64'h0000000000000000;
        dcache[651] <= 64'h0000000000000000;
        dcache[652] <= 64'h0000000000000000;
        dcache[653] <= 64'h0000000000000000;
        dcache[654] <= 64'h0000000000000000;
        dcache[655] <= 64'h0000000000000000;
        dcache[656] <= 64'h0000000000000000;
        dcache[657] <= 64'h0000000000000000;
        dcache[658] <= 64'h0000000000000000;
        dcache[659] <= 64'h0000000000000000;
        dcache[660] <= 64'h0000000000000000;
        dcache[661] <= 64'h0000000000000000;
        dcache[662] <= 64'h0000000000000000;
        dcache[663] <= 64'h0000000000000000;
        dcache[664] <= 64'h0000000000000000;
        dcache[665] <= 64'h0000000000000000;
        dcache[666] <= 64'h0000000000000000;
        dcache[667] <= 64'h0000000000000000;
        dcache[668] <= 64'h0000000000000000;
        dcache[669] <= 64'h0000000000000000;
        dcache[670] <= 64'h0000000000000000;
        dcache[671] <= 64'h0000000000000000;
        dcache[672] <= 64'h0000000000000000;
        dcache[673] <= 64'h0000000000000000;
        dcache[674] <= 64'h0000000000000000;
        dcache[675] <= 64'h0000000000000000;
        dcache[676] <= 64'h0000000000000000;
        dcache[677] <= 64'h0000000000000000;
        dcache[678] <= 64'h0000000000000000;
        dcache[679] <= 64'h0000000000000000;
        dcache[680] <= 64'h0000000000000000;
        dcache[681] <= 64'h0000000000000000;
        dcache[682] <= 64'h0000000000000000;
        dcache[683] <= 64'h0000000000000000;
        dcache[684] <= 64'h0000000000000000;
        dcache[685] <= 64'h0000000000000000;
        dcache[686] <= 64'h0000000000000000;
        dcache[687] <= 64'h0000000000000000;
        dcache[688] <= 64'h0000000000000000;
        dcache[689] <= 64'h0000000000000000;
        dcache[690] <= 64'h0000000000000000;
        dcache[691] <= 64'h0000000000000000;
        dcache[692] <= 64'h0000000000000000;
        dcache[693] <= 64'h0000000000000000;
        dcache[694] <= 64'h0000000000000000;
        dcache[695] <= 64'h0000000000000000;
        dcache[696] <= 64'h0000000000000000;
        dcache[697] <= 64'h0000000000000000;
        dcache[698] <= 64'h0000000000000000;
        dcache[699] <= 64'h0000000000000000;
        dcache[700] <= 64'h0000000000000000;
        dcache[701] <= 64'h0000000000000000;
        dcache[702] <= 64'h0000000000000000;
        dcache[703] <= 64'h0000000000000000;
        dcache[704] <= 64'h0000000000000000;
        dcache[705] <= 64'h0000000000000000;
        dcache[706] <= 64'h0000000000000000;
        dcache[707] <= 64'h0000000000000000;
        dcache[708] <= 64'h0000000000000000;
        dcache[709] <= 64'h0000000000000000;
        dcache[710] <= 64'h0000000000000000;
        dcache[711] <= 64'h0000000000000000;
        dcache[712] <= 64'h0000000000000000;
        dcache[713] <= 64'h0000000000000000;
        dcache[714] <= 64'h0000000000000000;
        dcache[715] <= 64'h0000000000000000;
        dcache[716] <= 64'h0000000000000000;
        dcache[717] <= 64'h0000000000000000;
        dcache[718] <= 64'h0000000000000000;
        dcache[719] <= 64'h0000000000000000;
        dcache[720] <= 64'h0000000000000000;
        dcache[721] <= 64'h0000000000000000;
        dcache[722] <= 64'h0000000000000000;
        dcache[723] <= 64'h0000000000000000;
        dcache[724] <= 64'h0000000000000000;
        dcache[725] <= 64'h0000000000000000;
        dcache[726] <= 64'h0000000000000000;
        dcache[727] <= 64'h0000000000000000;
        dcache[728] <= 64'h0000000000000000;
        dcache[729] <= 64'h0000000000000000;
        dcache[730] <= 64'h0000000000000000;
        dcache[731] <= 64'h0000000000000000;
        dcache[732] <= 64'h0000000000000000;
        dcache[733] <= 64'h0000000000000000;
        dcache[734] <= 64'h0000000000000000;
        dcache[735] <= 64'h0000000000000000;
        dcache[736] <= 64'h0000000000000000;
        dcache[737] <= 64'h0000000000000000;
        dcache[738] <= 64'h0000000000000000;
        dcache[739] <= 64'h0000000000000000;
        dcache[740] <= 64'h0000000000000000;
        dcache[741] <= 64'h0000000000000000;
        dcache[742] <= 64'h0000000000000000;
        dcache[743] <= 64'h0000000000000000;
        dcache[744] <= 64'h0000000000000000;
        dcache[745] <= 64'h0000000000000000;
        dcache[746] <= 64'h0000000000000000;
        dcache[747] <= 64'h0000000000000000;
        dcache[748] <= 64'h0000000000000000;
        dcache[749] <= 64'h0000000000000000;
        dcache[750] <= 64'h0000000000000000;
        dcache[751] <= 64'h0000000000000000;
        dcache[752] <= 64'h0000000000000000;
        dcache[753] <= 64'h0000000000000000;
        dcache[754] <= 64'h0000000000000000;
        dcache[755] <= 64'h0000000000000000;
        dcache[756] <= 64'h0000000000000000;
        dcache[757] <= 64'h0000000000000000;
        dcache[758] <= 64'h0000000000000000;
        dcache[759] <= 64'h0000000000000000;
        dcache[760] <= 64'h0000000000000000;
        dcache[761] <= 64'h0000000000000000;
        dcache[762] <= 64'h0000000000000000;
        dcache[763] <= 64'h0000000000000000;
        dcache[764] <= 64'h0000000000000000;
        dcache[765] <= 64'h0000000000000000;
        dcache[766] <= 64'h0000000000000000;
        dcache[767] <= 64'h0000000000000000;
        dcache[768] <= 64'h0000000000000000;
        dcache[769] <= 64'h0000000000000000;
        dcache[770] <= 64'h0000000000000000;
        dcache[771] <= 64'h0000000000000000;
        dcache[772] <= 64'h0000000000000000;
        dcache[773] <= 64'h0000000000000000;
        dcache[774] <= 64'h0000000000000000;
        dcache[775] <= 64'h0000000000000000;
        dcache[776] <= 64'h0000000000000000;
        dcache[777] <= 64'h0000000000000000;
        dcache[778] <= 64'h0000000000000000;
        dcache[779] <= 64'h0000000000000000;
        dcache[780] <= 64'h0000000000000000;
        dcache[781] <= 64'h0000000000000000;
        dcache[782] <= 64'h0000000000000000;
        dcache[783] <= 64'h0000000000000000;
        dcache[784] <= 64'h0000000000000000;
        dcache[785] <= 64'h0000000000000000;
        dcache[786] <= 64'h0000000000000000;
        dcache[787] <= 64'h0000000000000000;
        dcache[788] <= 64'h0000000000000000;
        dcache[789] <= 64'h0000000000000000;
        dcache[790] <= 64'h0000000000000000;
        dcache[791] <= 64'h0000000000000000;
        dcache[792] <= 64'h0000000000000000;
        dcache[793] <= 64'h0000000000000000;
        dcache[794] <= 64'h0000000000000000;
        dcache[795] <= 64'h0000000000000000;
        dcache[796] <= 64'h0000000000000000;
        dcache[797] <= 64'h0000000000000000;
        dcache[798] <= 64'h0000000000000000;
        dcache[799] <= 64'h0000000000000000;
        dcache[800] <= 64'h0000000000000000;
        dcache[801] <= 64'h0000000000000000;
        dcache[802] <= 64'h0000000000000000;
        dcache[803] <= 64'h0000000000000000;
        dcache[804] <= 64'h0000000000000000;
        dcache[805] <= 64'h0000000000000000;
        dcache[806] <= 64'h0000000000000000;
        dcache[807] <= 64'h0000000000000000;
        dcache[808] <= 64'h0000000000000000;
        dcache[809] <= 64'h0000000000000000;
        dcache[810] <= 64'h0000000000000000;
        dcache[811] <= 64'h0000000000000000;
        dcache[812] <= 64'h0000000000000000;
        dcache[813] <= 64'h0000000000000000;
        dcache[814] <= 64'h0000000000000000;
        dcache[815] <= 64'h0000000000000000;
        dcache[816] <= 64'h0000000000000000;
        dcache[817] <= 64'h0000000000000000;
        dcache[818] <= 64'h0000000000000000;
        dcache[819] <= 64'h0000000000000000;
        dcache[820] <= 64'h0000000000000000;
        dcache[821] <= 64'h0000000000000000;
        dcache[822] <= 64'h0000000000000000;
        dcache[823] <= 64'h0000000000000000;
        dcache[824] <= 64'h0000000000000000;
        dcache[825] <= 64'h0000000000000000;
        dcache[826] <= 64'h0000000000000000;
        dcache[827] <= 64'h0000000000000000;
        dcache[828] <= 64'h0000000000000000;
        dcache[829] <= 64'h0000000000000000;
        dcache[830] <= 64'h0000000000000000;
        dcache[831] <= 64'h0000000000000000;
        dcache[832] <= 64'h0000000000000000;
        dcache[833] <= 64'h0000000000000000;
        dcache[834] <= 64'h0000000000000000;
        dcache[835] <= 64'h0000000000000000;
        dcache[836] <= 64'h0000000000000000;
        dcache[837] <= 64'h0000000000000000;
        dcache[838] <= 64'h0000000000000000;
        dcache[839] <= 64'h0000000000000000;
        dcache[840] <= 64'h0000000000000000;
        dcache[841] <= 64'h0000000000000000;
        dcache[842] <= 64'h0000000000000000;
        dcache[843] <= 64'h0000000000000000;
        dcache[844] <= 64'h0000000000000000;
        dcache[845] <= 64'h0000000000000000;
        dcache[846] <= 64'h0000000000000000;
        dcache[847] <= 64'h0000000000000000;
        dcache[848] <= 64'h0000000000000000;
        dcache[849] <= 64'h0000000000000000;
        dcache[850] <= 64'h0000000000000000;
        dcache[851] <= 64'h0000000000000000;
        dcache[852] <= 64'h0000000000000000;
        dcache[853] <= 64'h0000000000000000;
        dcache[854] <= 64'h0000000000000000;
        dcache[855] <= 64'h0000000000000000;
        dcache[856] <= 64'h0000000000000000;
        dcache[857] <= 64'h0000000000000000;
        dcache[858] <= 64'h0000000000000000;
        dcache[859] <= 64'h0000000000000000;
        dcache[860] <= 64'h0000000000000000;
        dcache[861] <= 64'h0000000000000000;
        dcache[862] <= 64'h0000000000000000;
        dcache[863] <= 64'h0000000000000000;
        dcache[864] <= 64'h0000000000000000;
        dcache[865] <= 64'h0000000000000000;
        dcache[866] <= 64'h0000000000000000;
        dcache[867] <= 64'h0000000000000000;
        dcache[868] <= 64'h0000000000000000;
        dcache[869] <= 64'h0000000000000000;
        dcache[870] <= 64'h0000000000000000;
        dcache[871] <= 64'h0000000000000000;
        dcache[872] <= 64'h0000000000000000;
        dcache[873] <= 64'h0000000000000000;
        dcache[874] <= 64'h0000000000000000;
        dcache[875] <= 64'h0000000000000000;
        dcache[876] <= 64'h0000000000000000;
        dcache[877] <= 64'h0000000000000000;
        dcache[878] <= 64'h0000000000000000;
        dcache[879] <= 64'h0000000000000000;
        dcache[880] <= 64'h0000000000000000;
        dcache[881] <= 64'h0000000000000000;
        dcache[882] <= 64'h0000000000000000;
        dcache[883] <= 64'h0000000000000000;
        dcache[884] <= 64'h0000000000000000;
        dcache[885] <= 64'h0000000000000000;
        dcache[886] <= 64'h0000000000000000;
        dcache[887] <= 64'h0000000000000000;
        dcache[888] <= 64'h0000000000000000;
        dcache[889] <= 64'h0000000000000000;
        dcache[890] <= 64'h0000000000000000;
        dcache[891] <= 64'h0000000000000000;
        dcache[892] <= 64'h0000000000000000;
        dcache[893] <= 64'h0000000000000000;
        dcache[894] <= 64'h0000000000000000;
        dcache[895] <= 64'h0000000000000000;
        dcache[896] <= 64'h0000000000000000;
        dcache[897] <= 64'h0000000000000000;
        dcache[898] <= 64'h0000000000000000;
        dcache[899] <= 64'h0000000000000000;
        dcache[900] <= 64'h0000000000000000;
        dcache[901] <= 64'h0000000000000000;
        dcache[902] <= 64'h0000000000000000;
        dcache[903] <= 64'h0000000000000000;
        dcache[904] <= 64'h0000000000000000;
        dcache[905] <= 64'h0000000000000000;
        dcache[906] <= 64'h0000000000000000;
        dcache[907] <= 64'h0000000000000000;
        dcache[908] <= 64'h0000000000000000;
        dcache[909] <= 64'h0000000000000000;
        dcache[910] <= 64'h0000000000000000;
        dcache[911] <= 64'h0000000000000000;
        dcache[912] <= 64'h0000000000000000;
        dcache[913] <= 64'h0000000000000000;
        dcache[914] <= 64'h0000000000000000;
        dcache[915] <= 64'h0000000000000000;
        dcache[916] <= 64'h0000000000000000;
        dcache[917] <= 64'h0000000000000000;
        dcache[918] <= 64'h0000000000000000;
        dcache[919] <= 64'h0000000000000000;
        dcache[920] <= 64'h0000000000000000;
        dcache[921] <= 64'h0000000000000000;
        dcache[922] <= 64'h0000000000000000;
        dcache[923] <= 64'h0000000000000000;
        dcache[924] <= 64'h0000000000000000;
        dcache[925] <= 64'h0000000000000000;
        dcache[926] <= 64'h0000000000000000;
        dcache[927] <= 64'h0000000000000000;
        dcache[928] <= 64'h0000000000000000;
        dcache[929] <= 64'h0000000000000000;
        dcache[930] <= 64'h0000000000000000;
        dcache[931] <= 64'h0000000000000000;
        dcache[932] <= 64'h0000000000000000;
        dcache[933] <= 64'h0000000000000000;
        dcache[934] <= 64'h0000000000000000;
        dcache[935] <= 64'h0000000000000000;
        dcache[936] <= 64'h0000000000000000;
        dcache[937] <= 64'h0000000000000000;
        dcache[938] <= 64'h0000000000000000;
        dcache[939] <= 64'h0000000000000000;
        dcache[940] <= 64'h0000000000000000;
        dcache[941] <= 64'h0000000000000000;
        dcache[942] <= 64'h0000000000000000;
        dcache[943] <= 64'h0000000000000000;
        dcache[944] <= 64'h0000000000000000;
        dcache[945] <= 64'h0000000000000000;
        dcache[946] <= 64'h0000000000000000;
        dcache[947] <= 64'h0000000000000000;
        dcache[948] <= 64'h0000000000000000;
        dcache[949] <= 64'h0000000000000000;
        dcache[950] <= 64'h0000000000000000;
        dcache[951] <= 64'h0000000000000000;
        dcache[952] <= 64'h0000000000000000;
        dcache[953] <= 64'h0000000000000000;
        dcache[954] <= 64'h0000000000000000;
        dcache[955] <= 64'h0000000000000000;
        dcache[956] <= 64'h0000000000000000;
        dcache[957] <= 64'h0000000000000000;
        dcache[958] <= 64'h0000000000000000;
        dcache[959] <= 64'h0000000000000000;
        dcache[960] <= 64'h0000000000000000;
        dcache[961] <= 64'h0000000000000000;
        dcache[962] <= 64'h0000000000000000;
        dcache[963] <= 64'h0000000000000000;
        dcache[964] <= 64'h0000000000000000;
        dcache[965] <= 64'h0000000000000000;
        dcache[966] <= 64'h0000000000000000;
        dcache[967] <= 64'h0000000000000000;
        dcache[968] <= 64'h0000000000000000;
        dcache[969] <= 64'h0000000000000000;
        dcache[970] <= 64'h0000000000000000;
        dcache[971] <= 64'h0000000000000000;
        dcache[972] <= 64'h0000000000000000;
        dcache[973] <= 64'h0000000000000000;
        dcache[974] <= 64'h0000000000000000;
        dcache[975] <= 64'h0000000000000000;
        dcache[976] <= 64'h0000000000000000;
        dcache[977] <= 64'h0000000000000000;
        dcache[978] <= 64'h0000000000000000;
        dcache[979] <= 64'h0000000000000000;
        dcache[980] <= 64'h0000000000000000;
        dcache[981] <= 64'h0000000000000000;
        dcache[982] <= 64'h0000000000000000;
        dcache[983] <= 64'h0000000000000000;
        dcache[984] <= 64'h0000000000000000;
        dcache[985] <= 64'h0000000000000000;
        dcache[986] <= 64'h0000000000000000;
        dcache[987] <= 64'h0000000000000000;
        dcache[988] <= 64'h0000000000000000;
        dcache[989] <= 64'h0000000000000000;
        dcache[990] <= 64'h0000000000000000;
        dcache[991] <= 64'h0000000000000000;
        dcache[992] <= 64'h0000000000000000;
        dcache[993] <= 64'h0000000000000000;
        dcache[994] <= 64'h0000000000000000;
        dcache[995] <= 64'h0000000000000000;
        dcache[996] <= 64'h0000000000000000;
        dcache[997] <= 64'h0000000000000000;
        dcache[998] <= 64'h0000000000000000;
        dcache[999] <= 64'h0000000000000000;
        dcache[1000] <= 64'h0000000000000000;
        dcache[1001] <= 64'h0000000000000000;
        dcache[1002] <= 64'h0000000000000000;
        dcache[1003] <= 64'h0000000000000000;
        dcache[1004] <= 64'h0000000000000000;
        dcache[1005] <= 64'h0000000000000000;
        dcache[1006] <= 64'h0000000000000000;
        dcache[1007] <= 64'h0000000000000000;
        dcache[1008] <= 64'h0000000000000000;
        dcache[1009] <= 64'h0000000000000000;
        dcache[1010] <= 64'h0000000000000000;
        dcache[1011] <= 64'h0000000000000000;
        dcache[1012] <= 64'h0000000000000000;
        dcache[1013] <= 64'h0000000000000000;
        dcache[1014] <= 64'h0000000000000000;
        dcache[1015] <= 64'h0000000000000000;
        dcache[1016] <= 64'h0000000000000000;
        dcache[1017] <= 64'h0000000000000000;
        dcache[1018] <= 64'h0000000000000000;
        dcache[1019] <= 64'h0000000000000000;
        dcache[1020] <= 64'h0000000000000000;
        dcache[1021] <= 64'h0000000000000000;
        dcache[1022] <= 64'h0000000000000000;
        dcache[1023] <= 64'h0000000000000000;
    end

    initial begin
        $dumpfile("main_tb.vcd");
        $dumpvars(0, dcache[0]);
        $dumpvars(0, dcache[1]);
        $dumpvars(0, dcache[2]);
        $dumpvars(0, dcache[3]);
        $dumpvars(0, dcache[4]);
        $dumpvars(0, dcache[5]);
        $dumpvars(0, dcache[6]);
        $dumpvars(0, dcache[7]);
        $dumpvars(0, dcache[8]);
        $dumpvars(0, dcache[9]);
        $dumpvars(0, dcache[10]);
        $dumpvars(0, dcache[11]);
        $dumpvars(0, dcache[12]);
        $dumpvars(0, dcache[13]);
        $dumpvars(0, dcache[14]);
        $dumpvars(0, dcache[15]);
        $dumpvars(0, dcache[16]);
        $dumpvars(0, dcache[17]);
        $dumpvars(0, dcache[18]);
        $dumpvars(0, dcache[19]);
        $dumpvars(0, dcache[20]);
        $dumpvars(0, dcache[21]);
        $dumpvars(0, dcache[22]);
        $dumpvars(0, dcache[23]);
        $dumpvars(0, dcache[24]);
        $dumpvars(0, dcache[25]);
        $dumpvars(0, dcache[26]);
        $dumpvars(0, dcache[27]);
        $dumpvars(0, dcache[28]);
        $dumpvars(0, dcache[29]);
        $dumpvars(0, dcache[30]);
        $dumpvars(0, dcache[31]);
        $dumpvars(0, dcache[32]);
        $dumpvars(0, dcache[33]);
        $dumpvars(0, dcache[34]);
        $dumpvars(0, dcache[35]);
        $dumpvars(0, dcache[36]);
        $dumpvars(0, dcache[37]);
        $dumpvars(0, dcache[38]);
        $dumpvars(0, dcache[39]);
        $dumpvars(0, dcache[40]);
        $dumpvars(0, dcache[41]);
        $dumpvars(0, dcache[42]);
        $dumpvars(0, dcache[43]);
        $dumpvars(0, dcache[44]);
        $dumpvars(0, dcache[45]);
        $dumpvars(0, dcache[46]);
        $dumpvars(0, dcache[47]);
        $dumpvars(0, dcache[48]);
        $dumpvars(0, dcache[49]);
        $dumpvars(0, dcache[50]);
        $dumpvars(0, dcache[51]);
        $dumpvars(0, dcache[52]);
        $dumpvars(0, dcache[53]);
        $dumpvars(0, dcache[54]);
        $dumpvars(0, dcache[55]);
        $dumpvars(0, dcache[56]);
        $dumpvars(0, dcache[57]);
        $dumpvars(0, dcache[58]);
        $dumpvars(0, dcache[59]);
        $dumpvars(0, dcache[60]);
        $dumpvars(0, dcache[61]);
        $dumpvars(0, dcache[62]);
        $dumpvars(0, dcache[63]);
        $dumpvars(0, dcache[64]);
        $dumpvars(0, dcache[65]);
        $dumpvars(0, dcache[66]);
        $dumpvars(0, dcache[67]);
        $dumpvars(0, dcache[68]);
        $dumpvars(0, dcache[69]);
        $dumpvars(0, dcache[70]);
        $dumpvars(0, dcache[71]);
        $dumpvars(0, dcache[72]);
        $dumpvars(0, dcache[73]);
        $dumpvars(0, dcache[74]);
        $dumpvars(0, dcache[75]);
        $dumpvars(0, dcache[76]);
        $dumpvars(0, dcache[77]);
        $dumpvars(0, dcache[78]);
        $dumpvars(0, dcache[79]);
        $dumpvars(0, dcache[80]);
        $dumpvars(0, dcache[81]);
        $dumpvars(0, dcache[82]);
        $dumpvars(0, dcache[83]);
        $dumpvars(0, dcache[84]);
        $dumpvars(0, dcache[85]);
        $dumpvars(0, dcache[86]);
        $dumpvars(0, dcache[87]);
        $dumpvars(0, dcache[88]);
        $dumpvars(0, dcache[89]);
        $dumpvars(0, dcache[90]);
        $dumpvars(0, dcache[91]);
        $dumpvars(0, dcache[92]);
        $dumpvars(0, dcache[93]);
        $dumpvars(0, dcache[94]);
        $dumpvars(0, dcache[95]);
        $dumpvars(0, dcache[96]);
        $dumpvars(0, dcache[97]);
        $dumpvars(0, dcache[98]);
        $dumpvars(0, dcache[99]);
        $dumpvars(0, dcache[100]);
        $dumpvars(0, dcache[101]);
        $dumpvars(0, dcache[102]);
        $dumpvars(0, dcache[103]);
        $dumpvars(0, dcache[104]);
        $dumpvars(0, dcache[105]);
        $dumpvars(0, dcache[106]);
        $dumpvars(0, dcache[107]);
        $dumpvars(0, dcache[108]);
        $dumpvars(0, dcache[109]);
        $dumpvars(0, dcache[110]);
        $dumpvars(0, dcache[111]);
        $dumpvars(0, dcache[112]);
        $dumpvars(0, dcache[113]);
        $dumpvars(0, dcache[114]);
        $dumpvars(0, dcache[115]);
        $dumpvars(0, dcache[116]);
        $dumpvars(0, dcache[117]);
        $dumpvars(0, dcache[118]);
        $dumpvars(0, dcache[119]);
        $dumpvars(0, dcache[120]);
        $dumpvars(0, dcache[121]);
        $dumpvars(0, dcache[122]);
        $dumpvars(0, dcache[123]);
        $dumpvars(0, dcache[124]);
        $dumpvars(0, dcache[125]);
        $dumpvars(0, dcache[126]);
        $dumpvars(0, dcache[127]);
    end

endmodule
