module dcache_weights(address, read, data_out, valid, CLK, RST);
    parameter WIDTH = 32;
    parameter VEC_WIDTH = 64;
    reg [VEC_WIDTH-1:0] dcache [3191:0];
    
    input wire [WIDTH-1:0] address;
    input wire read;
    output wire [VEC_WIDTH-1:0] data_out;
    output wire valid;
    input CLK, RST;
    
    assign valid = 1'b1;
    
    wire [11:0] index = address[14:3];
    
    //always do this no matter what (read always active basically)
    assign data_out = dcache[index];
    
    initial begin
        dcache[0] = 64'h804b000b800c8013;
        dcache[1] = 64'h8007003700410000;
        dcache[2] = 64'h80158028803d8052;
        dcache[3] = 64'h00418024002a8026;
        dcache[4] = 64'h0014802a001e0022;
        dcache[5] = 64'h8013804b00420005;
        dcache[6] = 64'h0047800c002f8024;
        dcache[7] = 64'h804e80170033803d;
        dcache[8] = 64'h8001800f800a004a;
        dcache[9] = 64'h801c000100120030;
        dcache[10] = 64'h8045800f80228008;
        dcache[11] = 64'h800f001180100001;
        dcache[12] = 64'h802780578005004e;
        dcache[13] = 64'h002900510011002e;
        dcache[14] = 64'h003b803e80068035;
        dcache[15] = 64'h001b0048804e803d;
        dcache[16] = 64'h002300418058803b;
        dcache[17] = 64'h804a00440046001e;
        dcache[18] = 64'h005800450045003b;
        dcache[19] = 64'h0051805680538058;
        dcache[20] = 64'h00000020804e800a;
        dcache[21] = 64'h00520038800d803a;
        dcache[22] = 64'h000a80328038801b;
        dcache[23] = 64'h004400418025004f;
        dcache[24] = 64'h000d001f80530051;
        dcache[25] = 64'h0016804480120050;
        dcache[26] = 64'h003b000b803f0055;
        dcache[27] = 64'h8040004700480056;
        dcache[28] = 64'h8043003580250011;
        dcache[29] = 64'h8028001c80068054;
        dcache[30] = 64'h801d800e00518000;
        dcache[31] = 64'h8019004480358026;
        dcache[32] = 64'h80460037800c001a;
        dcache[33] = 64'h803180268015004c;
        dcache[34] = 64'h8011003b80190052;
        dcache[35] = 64'h0024801300508042;
        dcache[36] = 64'h004180288032004c;
        dcache[37] = 64'h8006000a0052801f;
        dcache[38] = 64'h0020804d000d0023;
        dcache[39] = 64'h8041004580450025;
        dcache[40] = 64'h8016804500040046;
        dcache[41] = 64'h8011804d804b804d;
        dcache[42] = 64'h803100508028800a;
        dcache[43] = 64'h8053003480430037;
        dcache[44] = 64'h8025800000558027;
        dcache[45] = 64'h001e800d80030033;
        dcache[46] = 64'h804d00488022802b;
        dcache[47] = 64'h003d800f00300012;
        dcache[48] = 64'h8016802980cf009c;
        dcache[49] = 64'h808c008a809180a8;
        dcache[50] = 64'h008200f4006c0086;
        dcache[51] = 64'h809780758080804f;
        dcache[52] = 64'h802600258075003a;
        dcache[53] = 64'h80e70064805e8054;
        dcache[54] = 64'h00fe00ea00820056;
        dcache[55] = 64'h80ff808980d6804f;
        dcache[56] = 64'h006480120015006c;
        dcache[57] = 64'h000f005e003300b4;
        dcache[58] = 64'h0026804780148093;
        dcache[59] = 64'h0052802e800f0024;
        dcache[60] = 64'h00278029004b803f;
        dcache[61] = 64'h006700058021802a;
        dcache[62] = 64'h004a8033800d001d;
        dcache[63] = 64'h0009002a00288024;
        dcache[64] = 64'h00458009004a803d;
        dcache[65] = 64'h80238044004a8058;
        dcache[66] = 64'h8054801400198055;
        dcache[67] = 64'h80138007002c0021;
        dcache[68] = 64'h0028800e00478037;
        dcache[69] = 64'h001c000f8030001d;
        dcache[70] = 64'h8045802e00048022;
        dcache[71] = 64'h003e803d00438006;
        dcache[72] = 64'h803e0055000d0051;
        dcache[73] = 64'h001a0045803a0026;
        dcache[74] = 64'h803b80490026804b;
        dcache[75] = 64'h0054003d8022804b;
        dcache[76] = 64'h0017804180008001;
        dcache[77] = 64'h803f800f80168009;
        dcache[78] = 64'h801e801a001f802d;
        dcache[79] = 64'h002c800100008009;
        dcache[80] = 64'h80178024801f0013;
        dcache[81] = 64'h000e805880468009;
        dcache[82] = 64'h00478035801b8010;
        dcache[83] = 64'h00328047000f8047;
        dcache[84] = 64'h004780270028800e;
        dcache[85] = 64'h8034805280398048;
        dcache[86] = 64'h8007004a8048801e;
        dcache[87] = 64'h00548019803c0048;
        dcache[88] = 64'h001f0018801b801b;
        dcache[89] = 64'h000e003b803b804d;
        dcache[90] = 64'h00488032003c0017;
        dcache[91] = 64'h8055002e8038801f;
        dcache[92] = 64'h000f0030004b8049;
        dcache[93] = 64'h8018800680468005;
        dcache[94] = 64'h80288037804c0033;
        dcache[95] = 64'h0010805700468010;
        dcache[96] = 64'h0056004980450017;
        dcache[97] = 64'h801100530045801c;
        dcache[98] = 64'h0034005700338009;
        dcache[99] = 64'h802c804d80348057;
        dcache[100] = 64'h0021004300330037;
        dcache[101] = 64'h003b801b00500011;
        dcache[102] = 64'h0021804400260007;
        dcache[103] = 64'h804d802180320024;
        dcache[104] = 64'h003500090016801c;
        dcache[105] = 64'h0011003380198030;
        dcache[106] = 64'h0049801a0002802b;
        dcache[107] = 64'h801b0003001a804a;
        dcache[108] = 64'h003b000e0027802a;
        dcache[109] = 64'h00218009804a0012;
        dcache[110] = 64'h000380260004004c;
        dcache[111] = 64'h0048800d002f0002;
        dcache[112] = 64'h8018801800248045;
        dcache[113] = 64'h803e000580128016;
        dcache[114] = 64'h80290015001f802a;
        dcache[115] = 64'h001a801e802e0041;
        dcache[116] = 64'h80110013804d8028;
        dcache[117] = 64'h804d002800050047;
        dcache[118] = 64'h8024004680328042;
        dcache[119] = 64'h0007004c00498012;
        dcache[120] = 64'h804a800400018052;
        dcache[121] = 64'h8028002c8018001c;
        dcache[122] = 64'h004b001880190051;
        dcache[123] = 64'h805480020039003b;
        dcache[124] = 64'h8056804b800c804d;
        dcache[125] = 64'h000f00040020803c;
        dcache[126] = 64'h800a0044000f8028;
        dcache[127] = 64'h0028001080318013;
        dcache[128] = 64'h80450055802f0060;
        dcache[129] = 64'h801a00808044002e;
        dcache[130] = 64'h0068009f005900b5;
        dcache[131] = 64'h8067801880498050;
        dcache[132] = 64'h8091004880c80050;
        dcache[133] = 64'h8094002b8047002e;
        dcache[134] = 64'h008b00c4006100a0;
        dcache[135] = 64'h8096805e80308025;
        dcache[136] = 64'h810680a7804e0143;
        dcache[137] = 64'h817100c3808a8061;
        dcache[138] = 64'h016900e80113017f;
        dcache[139] = 64'h819d804780c0802d;
        dcache[140] = 64'h8154808a80790165;
        dcache[141] = 64'h812d018680b3805d;
        dcache[142] = 64'h0172013a0114020b;
        dcache[143] = 64'h81b1000380d80004;
        dcache[144] = 64'h80c780bc8149016e;
        dcache[145] = 64'h818101258098803e;
        dcache[146] = 64'h01690168014b017f;
        dcache[147] = 64'h8136804180cd0055;
        dcache[148] = 64'h80d180ed816d0124;
        dcache[149] = 64'h81e401cd81098044;
        dcache[150] = 64'h023a01fc01640172;
        dcache[151] = 64'h81b7805c81040098;
        dcache[152] = 64'h8097815d81ca010d;
        dcache[153] = 64'h811202a080f0817f;
        dcache[154] = 64'h029c0235024a02cf;
        dcache[155] = 64'h82bf8039809500cf;
        dcache[156] = 64'h806d807f81a700e6;
        dcache[157] = 64'h8156008c80ee81a7;
        dcache[158] = 64'h020902670277021a;
        dcache[159] = 64'h812a0096810200d7;
        dcache[160] = 64'h8119812a81be0168;
        dcache[161] = 64'h81d30093810a816b;
        dcache[162] = 64'h02a5030d02a401e7;
        dcache[163] = 64'h8111003280d50082;
        dcache[164] = 64'h810480c381d30346;
        dcache[165] = 64'h81838034809681b4;
        dcache[166] = 64'h026000fd033302dd;
        dcache[167] = 64'h80ef0048812100f0;
        dcache[168] = 64'h804280e9006402d0;
        dcache[169] = 64'h8038806780fa80ec;
        dcache[170] = 64'h80f4804f01390187;
        dcache[171] = 64'h81ad012100760089;
        dcache[172] = 64'h813e81b200160280;
        dcache[173] = 64'h81ae802180f8000c;
        dcache[174] = 64'h008a020a018f00d8;
        dcache[175] = 64'h80f500d9808100cd;
        dcache[176] = 64'h81b6819680540294;
        dcache[177] = 64'h8136002f80260052;
        dcache[178] = 64'h0220015d013e0046;
        dcache[179] = 64'h805381058082007a;
        dcache[180] = 64'h813480a781310272;
        dcache[181] = 64'h811200b380318017;
        dcache[182] = 64'h0276024801fa00b8;
        dcache[183] = 64'h80de81a2812e8000;
        dcache[184] = 64'h810b8123816f01e2;
        dcache[185] = 64'h81a302e9810380ef;
        dcache[186] = 64'h01b3021701d6018f;
        dcache[187] = 64'h81de8174817d0075;
        dcache[188] = 64'h8145811281c200df;
        dcache[189] = 64'h817201ba814b80ff;
        dcache[190] = 64'h01d801b001a801f1;
        dcache[191] = 64'h81d8810b81040020;
        dcache[192] = 64'h8104810f812e005e;
        dcache[193] = 64'h817001218101814f;
        dcache[194] = 64'h0137017d015101be;
        dcache[195] = 64'h817f810a81098021;
        dcache[196] = 64'h80aa80e380c600c2;
        dcache[197] = 64'h811201ac80ba80f3;
        dcache[198] = 64'h0128010c00ae01b6;
        dcache[199] = 64'h817780d2815d801c;
        dcache[200] = 64'h80ce803b809f010b;
        dcache[201] = 64'h8105015280ba80ce;
        dcache[202] = 64'h00eb012600c70173;
        dcache[203] = 64'h8124807181678016;
        dcache[204] = 64'h8049805a802700f3;
        dcache[205] = 64'h808c00a880a40015;
        dcache[206] = 64'h013100d400b300e0;
        dcache[207] = 64'h8134805680d70018;
        dcache[208] = 64'h002e005480480054;
        dcache[209] = 64'h00350050001d004c;
        dcache[210] = 64'h0043801d80018005;
        dcache[211] = 64'h80138001001e803e;
        dcache[212] = 64'h0014004e00130024;
        dcache[213] = 64'h003680330005004c;
        dcache[214] = 64'h802e0046802b8030;
        dcache[215] = 64'h00258008801d0029;
        dcache[216] = 64'h00000050001d8010;
        dcache[217] = 64'h0017003e00550024;
        dcache[218] = 64'h802e80248056001c;
        dcache[219] = 64'h00018003003f8039;
        dcache[220] = 64'h001d803d0054802c;
        dcache[221] = 64'h001d001280238049;
        dcache[222] = 64'h8019803880410008;
        dcache[223] = 64'h80390038804f8057;
        dcache[224] = 64'h801b802000350028;
        dcache[225] = 64'h000c000800488027;
        dcache[226] = 64'h0055805080318054;
        dcache[227] = 64'h0001000c80290003;
        dcache[228] = 64'h8054003d0017003a;
        dcache[229] = 64'h8023805780260028;
        dcache[230] = 64'h0027002a00140040;
        dcache[231] = 64'h0014001000458006;
        dcache[232] = 64'h0009004d80c600f7;
        dcache[233] = 64'h808300628036802d;
        dcache[234] = 64'h006c006e004d801d;
        dcache[235] = 64'h80288023807e002c;
        dcache[236] = 64'h80dc806e80530033;
        dcache[237] = 64'h80b6810a00348024;
        dcache[238] = 64'h0133014c00a680c7;
        dcache[239] = 64'h008b007d80d38022;
        dcache[240] = 64'h8135810580e900e0;
        dcache[241] = 64'h814a80ba801a8095;
        dcache[242] = 64'h015a01d801268006;
        dcache[243] = 64'h0080008381088023;
        dcache[244] = 64'h80a480f5815d0107;
        dcache[245] = 64'h002601a800138032;
        dcache[246] = 64'h013b015801550147;
        dcache[247] = 64'h822b80dd80d30062;
        dcache[248] = 64'h815f807581820178;
        dcache[249] = 64'h0072012200128079;
        dcache[250] = 64'h024201a201d30104;
        dcache[251] = 64'h813000b781160074;
        dcache[252] = 64'h817d815981f5024c;
        dcache[253] = 64'h80c2027d00068022;
        dcache[254] = 64'h025c02c2028301f5;
        dcache[255] = 64'h8274802b81800018;
        dcache[256] = 64'h81cd801d818001e9;
        dcache[257] = 64'h804902f800ab80d0;
        dcache[258] = 64'h028301a3024d012b;
        dcache[259] = 64'h81ba80eb814e0025;
        dcache[260] = 64'h82c2007f81050133;
        dcache[261] = 64'h00d5048c01fb0075;
        dcache[262] = 64'h0177002901c2806f;
        dcache[263] = 64'h802981a1814e016c;
        dcache[264] = 64'h82dc8023809400a0;
        dcache[265] = 64'h000c04f002028068;
        dcache[266] = 64'h024d018802de005e;
        dcache[267] = 64'h809b826f81ff0168;
        dcache[268] = 64'h824780c4001f00da;
        dcache[269] = 64'h80300563021d0093;
        dcache[270] = 64'h015601f903f40165;
        dcache[271] = 64'h805681e682b30130;
        dcache[272] = 64'h822e8061005700c4;
        dcache[273] = 64'h801103de01b00098;
        dcache[274] = 64'h00df01a0037e011a;
        dcache[275] = 64'h80918133838a016b;
        dcache[276] = 64'h829b81b500490168;
        dcache[277] = 64'h809901c0008200fc;
        dcache[278] = 64'h80a2012302cd007d;
        dcache[279] = 64'h81d3001b82d10139;
        dcache[280] = 64'h829d81b10104016d;
        dcache[281] = 64'h802102ce012b00da;
        dcache[282] = 64'h800500ec04430103;
        dcache[283] = 64'h826081d5829d000d;
        dcache[284] = 64'h81b681d0025501f2;
        dcache[285] = 64'h804a033e00dc015b;
        dcache[286] = 64'h802b00bd0288001a;
        dcache[287] = 64'h8297810f82ce0019;
        dcache[288] = 64'h81af811c012802e1;
        dcache[289] = 64'h8044014f002e01a2;
        dcache[290] = 64'h809a00c500a40027;
        dcache[291] = 64'h814880b5829c0038;
        dcache[292] = 64'h80688123800402a1;
        dcache[293] = 64'h0085017980030083;
        dcache[294] = 64'h002201090066004e;
        dcache[295] = 64'h81f480b080be808b;
        dcache[296] = 64'h82598016001101f5;
        dcache[297] = 64'h00b200ce80660071;
        dcache[298] = 64'h00ab00f500778025;
        dcache[299] = 64'h81f0000700760008;
        dcache[300] = 64'h8239814781070324;
        dcache[301] = 64'h80440149804c805e;
        dcache[302] = 64'h803301f800a3012d;
        dcache[303] = 64'h81e2801500098003;
        dcache[304] = 64'h81cb80f881a601c4;
        dcache[305] = 64'h80c901bf003b804d;
        dcache[306] = 64'h003101f200fe015f;
        dcache[307] = 64'h82a480cd00180001;
        dcache[308] = 64'h809f813681f40013;
        dcache[309] = 64'h800601b60150803b;
        dcache[310] = 64'h01bb016502170147;
        dcache[311] = 64'h8263826c81540034;
        dcache[312] = 64'h003280fe822d00eb;
        dcache[313] = 64'h80ec0108008d81ba;
        dcache[314] = 64'h01d9015402800303;
        dcache[315] = 64'h81d782ab8181809b;
        dcache[316] = 64'h81a1000980570193;
        dcache[317] = 64'h810501df006e806d;
        dcache[318] = 64'h01730219020b803e;
        dcache[319] = 64'h80c382a9823d8007;
        dcache[320] = 64'h80aa0031009f000e;
        dcache[321] = 64'h00c001c00154802a;
        dcache[322] = 64'h0071805600a980c5;
        dcache[323] = 64'h00f081b7000b009f;
        dcache[324] = 64'h805a006a00b78054;
        dcache[325] = 64'h00c300d9013a0006;
        dcache[326] = 64'h807080f0009c8102;
        dcache[327] = 64'h011380dd0026006c;
        dcache[328] = 64'h8024003f803f8056;
        dcache[329] = 64'h8028804d00260024;
        dcache[330] = 64'h802b000d80420055;
        dcache[331] = 64'h001d804f00170003;
        dcache[332] = 64'h0041004c0011800b;
        dcache[333] = 64'h002e00478009004c;
        dcache[334] = 64'h8057002480150037;
        dcache[335] = 64'h800380130055802d;
        dcache[336] = 64'h8029804400568015;
        dcache[337] = 64'h00020056003f8018;
        dcache[338] = 64'h804c802c00140011;
        dcache[339] = 64'h804c800c801d8041;
        dcache[340] = 64'h0048800980020043;
        dcache[341] = 64'h000e000700060042;
        dcache[342] = 64'h803d0014001e802c;
        dcache[343] = 64'h8024803c8010804a;
        dcache[344] = 64'h001f808f005f0095;
        dcache[345] = 64'h8178004480570157;
        dcache[346] = 64'h80b20116009680e6;
        dcache[347] = 64'h80cc0117814280e5;
        dcache[348] = 64'h80fd80a28054007d;
        dcache[349] = 64'h81008055000000e6;
        dcache[350] = 64'h00c30159007c80f1;
        dcache[351] = 64'h0093007f80c1007c;
        dcache[352] = 64'h806e809881730018;
        dcache[353] = 64'h005b0001807a00fc;
        dcache[354] = 64'h801e021b00e40058;
        dcache[355] = 64'h802a003000120029;
        dcache[356] = 64'h8143009e00b481c6;
        dcache[357] = 64'h80ef005201010018;
        dcache[358] = 64'h808900f801d5018f;
        dcache[359] = 64'h019881978008807e;
        dcache[360] = 64'h823c013e00cc80c2;
        dcache[361] = 64'h003c01db019d0112;
        dcache[362] = 64'h8014018002040127;
        dcache[363] = 64'h8091814e8017811f;
        dcache[364] = 64'h831700e1009e808f;
        dcache[365] = 64'h00100198018901d2;
        dcache[366] = 64'h805e015500d401e7;
        dcache[367] = 64'h807f81558154808d;
        dcache[368] = 64'h83d0016a805f8117;
        dcache[369] = 64'h813f01be00dc016d;
        dcache[370] = 64'h002101b2006801a6;
        dcache[371] = 64'h0031820582150062;
        dcache[372] = 64'h83b800c000260077;
        dcache[373] = 64'h003a028901a80105;
        dcache[374] = 64'h00ec004200ab806f;
        dcache[375] = 64'h8043813982c800ef;
        dcache[376] = 64'h837f00e800ab80b8;
        dcache[377] = 64'h808001c600ea0087;
        dcache[378] = 64'h008b0065009800bd;
        dcache[379] = 64'h800d817d82390126;
        dcache[380] = 64'h830000b700758148;
        dcache[381] = 64'h806402390076009e;
        dcache[382] = 64'h012300e901430186;
        dcache[383] = 64'h009181e0829300fb;
        dcache[384] = 64'h840900c300e18010;
        dcache[385] = 64'h80bb021280230166;
        dcache[386] = 64'h808501bf0099012e;
        dcache[387] = 64'h001b815f825e019b;
        dcache[388] = 64'h84a9004700290122;
        dcache[389] = 64'h80640152808f00d6;
        dcache[390] = 64'h00cf013b01100086;
        dcache[391] = 64'h81108161821f02e3;
        dcache[392] = 64'h845600200023003d;
        dcache[393] = 64'h80d9008580b7005f;
        dcache[394] = 64'h008500a6004b012d;
        dcache[395] = 64'h804181f781520244;
        dcache[396] = 64'h838d004000950069;
        dcache[397] = 64'h80c4003d80c20079;
        dcache[398] = 64'h0049008c806000e1;
        dcache[399] = 64'h80b9813580b60129;
        dcache[400] = 64'h81fe814f009f8032;
        dcache[401] = 64'h80ed001a805f00ec;
        dcache[402] = 64'h003a006a80300067;
        dcache[403] = 64'h803681a980bb0116;
        dcache[404] = 64'h80ef80d200150047;
        dcache[405] = 64'h809580d080b200c6;
        dcache[406] = 64'h00e4005b80a2007b;
        dcache[407] = 64'h00c3815280080158;
        dcache[408] = 64'h813c80e7804a00c8;
        dcache[409] = 64'h80a28070810500a1;
        dcache[410] = 64'h005d011e80a70132;
        dcache[411] = 64'h80388149015a0147;
        dcache[412] = 64'h80c280c8802c022b;
        dcache[413] = 64'h80aa8031000500ce;
        dcache[414] = 64'h803a010f005a0130;
        dcache[415] = 64'h80bb81b9802700c4;
        dcache[416] = 64'h80730075804900c1;
        dcache[417] = 64'h8157809a00fd802e;
        dcache[418] = 64'h809d0182813c0190;
        dcache[419] = 64'h00298087809e0092;
        dcache[420] = 64'h804300e8811e0092;
        dcache[421] = 64'h80248080003f8132;
        dcache[422] = 64'h00ec014680d7012c;
        dcache[423] = 64'h817d805300568075;
        dcache[424] = 64'h8047009980d1007b;
        dcache[425] = 64'h01c2802580658206;
        dcache[426] = 64'h019300f38034007f;
        dcache[427] = 64'h822b00480101806a;
        dcache[428] = 64'h80bb007e80c6000b;
        dcache[429] = 64'h0012801780aa8373;
        dcache[430] = 64'h028501c500d8016d;
        dcache[431] = 64'h8154810700b580f6;
        dcache[432] = 64'h80e400ca80af00fe;
        dcache[433] = 64'h807900d0803681fd;
        dcache[434] = 64'h018b0194008b8045;
        dcache[435] = 64'h007c8163001400bb;
        dcache[436] = 64'h80020186801b00f8;
        dcache[437] = 64'h00d0003400758213;
        dcache[438] = 64'h8017802c80c3810d;
        dcache[439] = 64'h01a0005180310110;
        dcache[440] = 64'h0014003f80dd0117;
        dcache[441] = 64'h80090130011e812e;
        dcache[442] = 64'h007801000011011f;
        dcache[443] = 64'h00d0804380a800a3;
        dcache[444] = 64'h0035001c8007001f;
        dcache[445] = 64'h0044804c00248020;
        dcache[446] = 64'h8030804700338039;
        dcache[447] = 64'h0040802400140016;
        dcache[448] = 64'h0016800f8023801c;
        dcache[449] = 64'h80248009002d8006;
        dcache[450] = 64'h0036002d003f0014;
        dcache[451] = 64'h800700298057004c;
        dcache[452] = 64'h000c006a80288008;
        dcache[453] = 64'h80b980340001800f;
        dcache[454] = 64'h801d00808034006e;
        dcache[455] = 64'h0016000f800f8057;
        dcache[456] = 64'h0030003c019e80a9;
        dcache[457] = 64'h8182800480750111;
        dcache[458] = 64'h810a015900d58062;
        dcache[459] = 64'h00350074812c811b;
        dcache[460] = 64'h00fb013300f98189;
        dcache[461] = 64'h818580ca81bc00ad;
        dcache[462] = 64'h81e5019480e7016b;
        dcache[463] = 64'h019e806d00a00017;
        dcache[464] = 64'h8078800800e781b3;
        dcache[465] = 64'h809e00c600360003;
        dcache[466] = 64'h808e0136019401fc;
        dcache[467] = 64'h8009818800aa006c;
        dcache[468] = 64'h814c806201a880e5;
        dcache[469] = 64'h8050024000c40035;
        dcache[470] = 64'h8137010601e901f5;
        dcache[471] = 64'h8085820780a0808b;
        dcache[472] = 64'h824d010c01ca80ad;
        dcache[473] = 64'h00b2022a01880179;
        dcache[474] = 64'h80ac00c5004e009a;
        dcache[475] = 64'h804e8101801d0100;
        dcache[476] = 64'h82390169007d80b9;
        dcache[477] = 64'h00e000ff01190072;
        dcache[478] = 64'h008080c5803500ab;
        dcache[479] = 64'h801a808500970187;
        dcache[480] = 64'h829a009a01558020;
        dcache[481] = 64'h8027017e00f80043;
        dcache[482] = 64'h803100660158010f;
        dcache[483] = 64'h803281988102012f;
        dcache[484] = 64'h832c005201758075;
        dcache[485] = 64'h8017013a00978031;
        dcache[486] = 64'h005a804c00510054;
        dcache[487] = 64'h005d80fb815e0182;
        dcache[488] = 64'h82e9010701368092;
        dcache[489] = 64'h80890134001c807d;
        dcache[490] = 64'h800c008f002a0117;
        dcache[491] = 64'h803d809c813600de;
        dcache[492] = 64'h817c011500a48009;
        dcache[493] = 64'h0066003e000a800f;
        dcache[494] = 64'h000d001f80f50096;
        dcache[495] = 64'h0079803080590281;
        dcache[496] = 64'h810e009f013680a7;
        dcache[497] = 64'h008a0051006c8091;
        dcache[498] = 64'h80018080804e0096;
        dcache[499] = 64'h8059801780df01c0;
        dcache[500] = 64'h81b500560166801b;
        dcache[501] = 64'h801a003e00250008;
        dcache[502] = 64'h0021807480a200e1;
        dcache[503] = 64'h8046805381780179;
        dcache[504] = 64'h827e003e013d8015;
        dcache[505] = 64'h0005002e00340054;
        dcache[506] = 64'h005a802080720066;
        dcache[507] = 64'h80820059801e0195;
        dcache[508] = 64'h812d009500510036;
        dcache[509] = 64'h8073801b80498002;
        dcache[510] = 64'h001b8005818f00c2;
        dcache[511] = 64'h80530007801c01ba;
        dcache[512] = 64'h001600b100888031;
        dcache[513] = 64'h8087008f80e40050;
        dcache[514] = 64'h0068003e804d001e;
        dcache[515] = 64'h814080cb0002012a;
        dcache[516] = 64'h001200410068002a;
        dcache[517] = 64'h0072006180b6803d;
        dcache[518] = 64'h00a30024806e001d;
        dcache[519] = 64'h801e807d008b00c4;
        dcache[520] = 64'h8097008b003b008f;
        dcache[521] = 64'h00180043808b006b;
        dcache[522] = 64'h0089009180a58019;
        dcache[523] = 64'h00388014008b00e1;
        dcache[524] = 64'h010a006480368019;
        dcache[525] = 64'h004600bc802b00cb;
        dcache[526] = 64'h00620017000400b7;
        dcache[527] = 64'h8049804e00040023;
        dcache[528] = 64'h00bb0028805680ba;
        dcache[529] = 64'h800a007c002500d1;
        dcache[530] = 64'h00a8803080df009f;
        dcache[531] = 64'h8025804c8108803e;
        dcache[532] = 64'h0198006680eb006c;
        dcache[533] = 64'h00a4000480d0006a;
        dcache[534] = 64'h008d002780dc0181;
        dcache[535] = 64'h807c00d48040800b;
        dcache[536] = 64'h006e007a812b003d;
        dcache[537] = 64'h8008810e808a801f;
        dcache[538] = 64'h00c68029814f019a;
        dcache[539] = 64'h80710002007e80b2;
        dcache[540] = 64'h805e80098227800a;
        dcache[541] = 64'h8042807c0013815f;
        dcache[542] = 64'h00db004781030150;
        dcache[543] = 64'h80ff000700878181;
        dcache[544] = 64'h001c021c80d180c6;
        dcache[545] = 64'h031780f5008381da;
        dcache[546] = 64'h801180ab80fa00c9;
        dcache[547] = 64'h00140080018e8018;
        dcache[548] = 64'h804c027f008400ab;
        dcache[549] = 64'h01be80c58091820c;
        dcache[550] = 64'h00220026808d8043;
        dcache[551] = 64'h00c90055019c009e;
        dcache[552] = 64'h80ff00ca011c018a;
        dcache[553] = 64'h0079814081b781e4;
        dcache[554] = 64'h00be019400e380e8;
        dcache[555] = 64'h010c00ac01980138;
        dcache[556] = 64'h80b1804e80a90023;
        dcache[557] = 64'h001a00e4800e817e;
        dcache[558] = 64'h017c018001400065;
        dcache[559] = 64'h803e8179008d80c0;
        dcache[560] = 64'h003d004b00208036;
        dcache[561] = 64'h8056002480288016;
        dcache[562] = 64'h803f00538014801c;
        dcache[563] = 64'h8027800080450040;
        dcache[564] = 64'h8017001000560042;
        dcache[565] = 64'h8047002280270005;
        dcache[566] = 64'h0025003d00418031;
        dcache[567] = 64'h0010804a80278029;
        dcache[568] = 64'h805e80fc02130076;
        dcache[569] = 64'h811501ff812a0177;
        dcache[570] = 64'h802901de01260032;
        dcache[571] = 64'h811e80a581dd80b9;
        dcache[572] = 64'h0033007a021a811a;
        dcache[573] = 64'h803300db000f00c0;
        dcache[574] = 64'h810e004b00360049;
        dcache[575] = 64'h011100158111011f;
        dcache[576] = 64'h80c280b3021781ae;
        dcache[577] = 64'h809e021301890067;
        dcache[578] = 64'h806c002e02ff0114;
        dcache[579] = 64'h00cf8160803f0063;
        dcache[580] = 64'h005e00540154807e;
        dcache[581] = 64'h801d002f801f00ef;
        dcache[582] = 64'h826100e001630111;
        dcache[583] = 64'h00bd807c810780db;
        dcache[584] = 64'h814c007f00c980af;
        dcache[585] = 64'h8024805000fe0038;
        dcache[586] = 64'h8084007e00a00105;
        dcache[587] = 64'h0060805480ca0063;
        dcache[588] = 64'h811800ee00a780c7;
        dcache[589] = 64'h8016007500018086;
        dcache[590] = 64'h8074005e00b200b7;
        dcache[591] = 64'h000580b880bf00a4;
        dcache[592] = 64'h8027003c807f8086;
        dcache[593] = 64'h0079003300738064;
        dcache[594] = 64'h803980a3019000ee;
        dcache[595] = 64'h003681de804d0123;
        dcache[596] = 64'h008a00a90019806d;
        dcache[597] = 64'h0085008200b80012;
        dcache[598] = 64'h809680d8007600a4;
        dcache[599] = 64'h001c808880380018;
        dcache[600] = 64'h00028072809400bc;
        dcache[601] = 64'h00a88020001e8048;
        dcache[602] = 64'h002e8031801800c5;
        dcache[603] = 64'h001b80b68001011e;
        dcache[604] = 64'h806280b5006a8025;
        dcache[605] = 64'h00e5807b00000029;
        dcache[606] = 64'h004b80738003003a;
        dcache[607] = 64'h0110804f0177015a;
        dcache[608] = 64'h0009801100c80039;
        dcache[609] = 64'h0130804c80ac801f;
        dcache[610] = 64'h803e813a80000095;
        dcache[611] = 64'h00e9805e011b013f;
        dcache[612] = 64'h80b5801600a30017;
        dcache[613] = 64'h005c80ec80aa8063;
        dcache[614] = 64'h000200188039004e;
        dcache[615] = 64'h00ad006500150177;
        dcache[616] = 64'h8015001000ad0039;
        dcache[617] = 64'h8072000f806d8042;
        dcache[618] = 64'h00518032808b0078;
        dcache[619] = 64'h8001803900070112;
        dcache[620] = 64'h0019806a01060029;
        dcache[621] = 64'h8026803700250049;
        dcache[622] = 64'h0021804b80a00070;
        dcache[623] = 64'h8046805680d000de;
        dcache[624] = 64'h0061004700d58001;
        dcache[625] = 64'h8038002b802e0093;
        dcache[626] = 64'h00b4808781450034;
        dcache[627] = 64'h8062809d0001011b;
        dcache[628] = 64'h805d00500036006f;
        dcache[629] = 64'h003b804080d98049;
        dcache[630] = 64'h00ad805d80ec803b;
        dcache[631] = 64'h8088802c007100f3;
        dcache[632] = 64'h80468032803700c1;
        dcache[633] = 64'h000a803d8017801d;
        dcache[634] = 64'h008e804980f60074;
        dcache[635] = 64'h808180e6800f006e;
        dcache[636] = 64'h8022800c00760063;
        dcache[637] = 64'h0000002680738022;
        dcache[638] = 64'h003480068032010a;
        dcache[639] = 64'h8092803900720013;
        dcache[640] = 64'h80af00bc0047801a;
        dcache[641] = 64'h00568024809e0067;
        dcache[642] = 64'h008c00528112003c;
        dcache[643] = 64'h812e004a008f0087;
        dcache[644] = 64'h00250012002c800e;
        dcache[645] = 64'h00b0802380a6004a;
        dcache[646] = 64'h0063006a8083801f;
        dcache[647] = 64'h8135006180a6002d;
        dcache[648] = 64'h011c806c80b70032;
        dcache[649] = 64'h804400358095016e;
        dcache[650] = 64'h8007808f80bf0081;
        dcache[651] = 64'h80af0083807100b2;
        dcache[652] = 64'h0077808f817b8008;
        dcache[653] = 64'h8009014d00d200bc;
        dcache[654] = 64'h80d5800c00330158;
        dcache[655] = 64'h8107801181288070;
        dcache[656] = 64'h006b009880660019;
        dcache[657] = 64'h01b100fc00828095;
        dcache[658] = 64'h802900d500520138;
        dcache[659] = 64'h8026800080548060;
        dcache[660] = 64'h8056019e017f00b1;
        dcache[661] = 64'h0382801b004881a5;
        dcache[662] = 64'h0107006b004a002e;
        dcache[663] = 64'h801380d0013e01f9;
        dcache[664] = 64'h8074011080370076;
        dcache[665] = 64'h026b004080218184;
        dcache[666] = 64'h006f0185010300af;
        dcache[667] = 64'h8195807a0168804c;
        dcache[668] = 64'h00e8000c805a010f;
        dcache[669] = 64'h00c00197809580f8;
        dcache[670] = 64'h0105011800d500fc;
        dcache[671] = 64'h808980ad80718138;
        dcache[672] = 64'h000a003800310004;
        dcache[673] = 64'h8043801a00470043;
        dcache[674] = 64'h803f803180038044;
        dcache[675] = 64'h0046805180488058;
        dcache[676] = 64'h80a9007200d880cb;
        dcache[677] = 64'h80af006f809e00bd;
        dcache[678] = 64'h812e00f080e900d2;
        dcache[679] = 64'h010b80ab0020007e;
        dcache[680] = 64'h00bb014481760062;
        dcache[681] = 64'h8058000f80b70148;
        dcache[682] = 64'h00760078806200b2;
        dcache[683] = 64'h01cf801800cb006b;
        dcache[684] = 64'h012500cb00ee8262;
        dcache[685] = 64'h80ed001c00070038;
        dcache[686] = 64'h80c4001d018a8011;
        dcache[687] = 64'h01f080b681480154;
        dcache[688] = 64'h006c0084000080be;
        dcache[689] = 64'h001e020101030012;
        dcache[690] = 64'h800d8009012300c6;
        dcache[691] = 64'h8033806d00280072;
        dcache[692] = 64'h015300c580898072;
        dcache[693] = 64'h809a01ec80b80111;
        dcache[694] = 64'h8110804c807c00cc;
        dcache[695] = 64'h801180d48086800c;
        dcache[696] = 64'h005e00ae803580de;
        dcache[697] = 64'h80fc005f808d0103;
        dcache[698] = 64'h80cf8086003000dd;
        dcache[699] = 64'h012280ee80fc00ec;
        dcache[700] = 64'h0078002780528068;
        dcache[701] = 64'h0047804b80150070;
        dcache[702] = 64'h0042808401420059;
        dcache[703] = 64'h0075813680ba0064;
        dcache[704] = 64'h00d30034801a8049;
        dcache[705] = 64'h007f80a7805f8017;
        dcache[706] = 64'h808c802a00bf0090;
        dcache[707] = 64'h002e813b00670034;
        dcache[708] = 64'h00510107802f8044;
        dcache[709] = 64'h00838067807c0077;
        dcache[710] = 64'h80e5800300370082;
        dcache[711] = 64'h00d1811100fe8038;
        dcache[712] = 64'h8060007f001b005e;
        dcache[713] = 64'h007d805280b80171;
        dcache[714] = 64'h804b002680038058;
        dcache[715] = 64'h00a280ec005400e1;
        dcache[716] = 64'h801f806c002f0043;
        dcache[717] = 64'h005a8127803e0047;
        dcache[718] = 64'h000e00570028002a;
        dcache[719] = 64'h0128003e00390045;
        dcache[720] = 64'h807f0065006d00c8;
        dcache[721] = 64'h00f880bf80ab8024;
        dcache[722] = 64'h802f800e008c000f;
        dcache[723] = 64'h01410030004300a8;
        dcache[724] = 64'h80cf8056005b006c;
        dcache[725] = 64'h801280ee80240021;
        dcache[726] = 64'h0003002f80158020;
        dcache[727] = 64'h0152806100a200d1;
        dcache[728] = 64'h8079807b001f00d8;
        dcache[729] = 64'h00a1812f001f003b;
        dcache[730] = 64'h801c0093800d0064;
        dcache[731] = 64'h00f1802700c90157;
        dcache[732] = 64'h80cc804f002000a0;
        dcache[733] = 64'h00bd80e180390051;
        dcache[734] = 64'h000d00a800410013;
        dcache[735] = 64'h00c980e700c6017b;
        dcache[736] = 64'h8117806f00700018;
        dcache[737] = 64'h007180b8002f00aa;
        dcache[738] = 64'h0009005b0034006e;
        dcache[739] = 64'h00bb80f5004900f3;
        dcache[740] = 64'h8044805d00148035;
        dcache[741] = 64'h008d8166008d8048;
        dcache[742] = 64'h8034004400900022;
        dcache[743] = 64'h001c806a007400f4;
        dcache[744] = 64'h80fd802e00170054;
        dcache[745] = 64'h80018132002f000c;
        dcache[746] = 64'h8087008e80bc0002;
        dcache[747] = 64'h00bf800f000e00c9;
        dcache[748] = 64'h80a7004e802a0098;
        dcache[749] = 64'h007d811880ae0049;
        dcache[750] = 64'h002480ac80790029;
        dcache[751] = 64'h8012004800fd005a;
        dcache[752] = 64'h80ec00698018006f;
        dcache[753] = 64'h00158141807a004f;
        dcache[754] = 64'h8020801c80b80057;
        dcache[755] = 64'h802d00440076003f;
        dcache[756] = 64'h004b80278054801e;
        dcache[757] = 64'h807d8116008a802c;
        dcache[758] = 64'h0002807e008a801e;
        dcache[759] = 64'h007d001a807900aa;
        dcache[760] = 64'h00ec000380e8802b;
        dcache[761] = 64'h808d80398065004f;
        dcache[762] = 64'h005780ad8077004c;
        dcache[763] = 64'h800b00b100330149;
        dcache[764] = 64'h00d3800880368022;
        dcache[765] = 64'h8009004380ac802e;
        dcache[766] = 64'h007d80e80027015e;
        dcache[767] = 64'h80bd00e2000b0011;
        dcache[768] = 64'h002400fc8133015c;
        dcache[769] = 64'h013e01b380da80a4;
        dcache[770] = 64'h805a013380a50209;
        dcache[771] = 64'h814c003480270009;
        dcache[772] = 64'h808101a300d70244;
        dcache[773] = 64'h016300f8805c838b;
        dcache[774] = 64'h005b025c803f003b;
        dcache[775] = 64'h82720012020b00e6;
        dcache[776] = 64'h002c0129000901b6;
        dcache[777] = 64'h0160014c00c48211;
        dcache[778] = 64'h805100cb800900f2;
        dcache[779] = 64'h828a00ad0142003d;
        dcache[780] = 64'h014b802c806f013b;
        dcache[781] = 64'h8063012d00fd80fb;
        dcache[782] = 64'h003a014e007b00e7;
        dcache[783] = 64'h0002809d80958081;
        dcache[784] = 64'h8008802a80648003;
        dcache[785] = 64'h0035005200360030;
        dcache[786] = 64'h801b803a0027800b;
        dcache[787] = 64'h00198045806e0016;
        dcache[788] = 64'h802901600070012f;
        dcache[789] = 64'h8168013e81490150;
        dcache[790] = 64'h8177806780d80234;
        dcache[791] = 64'h014881fe00d00158;
        dcache[792] = 64'h00ee015b815180c3;
        dcache[793] = 64'h80000018809900f2;
        dcache[794] = 64'h0042807f806d0002;
        dcache[795] = 64'h01ef807100d50052;
        dcache[796] = 64'h02f400a50098823c;
        dcache[797] = 64'h80258055819500d2;
        dcache[798] = 64'h8088802d01ff803c;
        dcache[799] = 64'h0288810081580088;
        dcache[800] = 64'h008f0071026e81dc;
        dcache[801] = 64'h809103008001012b;
        dcache[802] = 64'h0066805d00ef005f;
        dcache[803] = 64'h004681648154016d;
        dcache[804] = 64'h003e00f6007b80aa;
        dcache[805] = 64'h80700180811d00cc;
        dcache[806] = 64'h80418206813d013c;
        dcache[807] = 64'h807180d3007b0094;
        dcache[808] = 64'h0064009d80178092;
        dcache[809] = 64'h0019804680b20058;
        dcache[810] = 64'h801e80df009c800b;
        dcache[811] = 64'h0112815d000e0072;
        dcache[812] = 64'h007700828065003e;
        dcache[813] = 64'h00240027813700a4;
        dcache[814] = 64'h804780b9009a0005;
        dcache[815] = 64'h800a80fb80608008;
        dcache[816] = 64'h0044010100220034;
        dcache[817] = 64'h0103807880df0133;
        dcache[818] = 64'h8023804e80878022;
        dcache[819] = 64'h8005816801a20020;
        dcache[820] = 64'h00c0008a803d8005;
        dcache[821] = 64'h001480a48048007c;
        dcache[822] = 64'h0035002e00600044;
        dcache[823] = 64'h007c80c400818017;
        dcache[824] = 64'h006300c180160077;
        dcache[825] = 64'h006580d780e000f9;
        dcache[826] = 64'h00c90057803d8040;
        dcache[827] = 64'h00c800e1008a008d;
        dcache[828] = 64'h8071004e806800ac;
        dcache[829] = 64'h00978081805c00d3;
        dcache[830] = 64'h0073003a802f8035;
        dcache[831] = 64'h01070068803f0099;
        dcache[832] = 64'h809f0064801f00ba;
        dcache[833] = 64'h000f80ee807e0079;
        dcache[834] = 64'h0038003a0054800e;
        dcache[835] = 64'h019d0067001f8012;
        dcache[836] = 64'h80ad8015005a00aa;
        dcache[837] = 64'h003d810880280102;
        dcache[838] = 64'h0037004e002f801a;
        dcache[839] = 64'h017d800200a1008c;
        dcache[840] = 64'h80e580b1801f019b;
        dcache[841] = 64'h0039803900430105;
        dcache[842] = 64'h804101150087004c;
        dcache[843] = 64'h014780260083011a;
        dcache[844] = 64'h804e80e1009a0057;
        dcache[845] = 64'h008a810900020017;
        dcache[846] = 64'h000300f900d000a3;
        dcache[847] = 64'h00dc805001380173;
        dcache[848] = 64'h803480ff003f00a1;
        dcache[849] = 64'h009d81c0002a0060;
        dcache[850] = 64'h808700a00001800b;
        dcache[851] = 64'h0046008d004f014a;
        dcache[852] = 64'h009480c4802c8031;
        dcache[853] = 64'h8018810d004900c6;
        dcache[854] = 64'h0008800880510071;
        dcache[855] = 64'h008c006e001600bb;
        dcache[856] = 64'h00c8801780520061;
        dcache[857] = 64'h808980fc00270018;
        dcache[858] = 64'h0033800e804c8038;
        dcache[859] = 64'h0042006500630152;
        dcache[860] = 64'h00610026002e0079;
        dcache[861] = 64'h009880eb80d70110;
        dcache[862] = 64'h8047807280b1804a;
        dcache[863] = 64'h004b006c8028010b;
        dcache[864] = 64'h800c804400670114;
        dcache[865] = 64'h003680f98042801f;
        dcache[866] = 64'h802f0011804d003c;
        dcache[867] = 64'h005100bc80160034;
        dcache[868] = 64'h001a806e80500074;
        dcache[869] = 64'h004c81020024802f;
        dcache[870] = 64'h00508058003e8070;
        dcache[871] = 64'h8076007900090073;
        dcache[872] = 64'h00f2005080980011;
        dcache[873] = 64'h00420008804a00e2;
        dcache[874] = 64'h0054808d806f8005;
        dcache[875] = 64'h80ae006a005a00d2;
        dcache[876] = 64'h00d3006680dd8018;
        dcache[877] = 64'h802a813a80ad807f;
        dcache[878] = 64'h00be80c6804d00b6;
        dcache[879] = 64'h80ae015a00d60040;
        dcache[880] = 64'h00fc00fc817b0160;
        dcache[881] = 64'h803b009380768152;
        dcache[882] = 64'h01088036814800b9;
        dcache[883] = 64'h80ee002e00af8066;
        dcache[884] = 64'h806900f700420157;
        dcache[885] = 64'h00bc0112002e8238;
        dcache[886] = 64'h00e701048151007c;
        dcache[887] = 64'h81b500b0021100c6;
        dcache[888] = 64'h01c7001200110136;
        dcache[889] = 64'h011d01b400e881cf;
        dcache[890] = 64'h808b80238017012d;
        dcache[891] = 64'h82ce00a0800d005b;
        dcache[892] = 64'h01470044819200a9;
        dcache[893] = 64'h002700cb010880fb;
        dcache[894] = 64'h006a019d80300129;
        dcache[895] = 64'h801c8036802180cc;
        dcache[896] = 64'h80c380f781080030;
        dcache[897] = 64'h812e0081006a0046;
        dcache[898] = 64'h011381448056814d;
        dcache[899] = 64'h00f700f080210002;
        dcache[900] = 64'h01ca01e281e9000c;
        dcache[901] = 64'h010e807f805e00cd;
        dcache[902] = 64'h8097002e01cd81a2;
        dcache[903] = 64'h024b81d781dc8000;
        dcache[904] = 64'h011800fa809e812b;
        dcache[905] = 64'h0090012e801400ae;
        dcache[906] = 64'h8004815380e8005c;
        dcache[907] = 64'h0054807700b2807d;
        dcache[908] = 64'h013400d7020e8216;
        dcache[909] = 64'h806600728166013a;
        dcache[910] = 64'h801280c8009a0086;
        dcache[911] = 64'h009e80f980360015;
        dcache[912] = 64'h0072007e02828174;
        dcache[913] = 64'h80760152820c0163;
        dcache[914] = 64'h801f80b001400095;
        dcache[915] = 64'h00068238811200b1;
        dcache[916] = 64'h00f500bf00c9809b;
        dcache[917] = 64'h0058801f81620073;
        dcache[918] = 64'h803480b800c7005c;
        dcache[919] = 64'h002580d500d18089;
        dcache[920] = 64'h00ba0078002a8041;
        dcache[921] = 64'h007e807980b680ca;
        dcache[922] = 64'h8027809e0105001c;
        dcache[923] = 64'h0059810a014c8084;
        dcache[924] = 64'h00a401380024800d;
        dcache[925] = 64'h0015802881e50050;
        dcache[926] = 64'h804a80cf011c806d;
        dcache[927] = 64'h004d812700958030;
        dcache[928] = 64'h010d009780d50021;
        dcache[929] = 64'h0035814b81440044;
        dcache[930] = 64'h0072004301498081;
        dcache[931] = 64'h00ab80ed00e68037;
        dcache[932] = 64'h00e700b5808c0062;
        dcache[933] = 64'h003a809080cd00a3;
        dcache[934] = 64'h0173805100718014;
        dcache[935] = 64'h80038003013e803e;
        dcache[936] = 64'h0080005a0035008a;
        dcache[937] = 64'h802d805680d700da;
        dcache[938] = 64'h00ba005a0050808a;
        dcache[939] = 64'h00c8002d00a98071;
        dcache[940] = 64'h0034011a80d1008f;
        dcache[941] = 64'h007c80c280c00169;
        dcache[942] = 64'h00e6001e80298017;
        dcache[943] = 64'h00bd00c5001c80d0;
        dcache[944] = 64'h800801298007007e;
        dcache[945] = 64'h0004809380b60080;
        dcache[946] = 64'h00e88028004b8068;
        dcache[947] = 64'h012e00cd80070040;
        dcache[948] = 64'h80a900e200b600b0;
        dcache[949] = 64'h803e80c200230090;
        dcache[950] = 64'h00ba800f00c5000f;
        dcache[951] = 64'h005300ce0005801d;
        dcache[952] = 64'h808b803a00450125;
        dcache[953] = 64'h808580c1802e0101;
        dcache[954] = 64'h8005006901128016;
        dcache[955] = 64'h011900850027010e;
        dcache[956] = 64'h802e801c003d0090;
        dcache[957] = 64'h803480b9805900f9;
        dcache[958] = 64'h802b802a00a78003;
        dcache[959] = 64'h01940028002900fe;
        dcache[960] = 64'h802280810031800c;
        dcache[961] = 64'h000680ec8015005c;
        dcache[962] = 64'h806e00078017804e;
        dcache[963] = 64'h0168001d00be0255;
        dcache[964] = 64'h000e80600047804a;
        dcache[965] = 64'h8009803e80670098;
        dcache[966] = 64'h8064000980938063;
        dcache[967] = 64'h00480067000901b3;
        dcache[968] = 64'h00d5002b0018809b;
        dcache[969] = 64'h806980c780900074;
        dcache[970] = 64'h001b806180298007;
        dcache[971] = 64'h011900fc00ca0135;
        dcache[972] = 64'h0048008200e88047;
        dcache[973] = 64'h804c8077804c008b;
        dcache[974] = 64'h8040806780b28070;
        dcache[975] = 64'h00800109004f00ef;
        dcache[976] = 64'h008c00e3807d801b;
        dcache[977] = 64'h80a700218051007f;
        dcache[978] = 64'h001e8055806e8038;
        dcache[979] = 64'h00490164004600f2;
        dcache[980] = 64'h004e009e8073801b;
        dcache[981] = 64'h808680cb80758085;
        dcache[982] = 64'h0002800080280001;
        dcache[983] = 64'h801f00bd002e0087;
        dcache[984] = 64'h001a00f280748046;
        dcache[985] = 64'h8099803180c000f6;
        dcache[986] = 64'h8004002800450029;
        dcache[987] = 64'h004900c200c70151;
        dcache[988] = 64'h017e0130821200d9;
        dcache[989] = 64'h807f803480e20056;
        dcache[990] = 64'h00c18150006d81a7;
        dcache[991] = 64'h001f01a200f70106;
        dcache[992] = 64'h018a015681848035;
        dcache[993] = 64'h0007814580668272;
        dcache[994] = 64'h00fc803880f7807b;
        dcache[995] = 64'h8123033f01df00b6;
        dcache[996] = 64'h00fc018c8021800a;
        dcache[997] = 64'h024600e580558211;
        dcache[998] = 64'h00898032806a0184;
        dcache[999] = 64'h830c033403b580ae;
        dcache[1000] = 64'h800902430165011f;
        dcache[1001] = 64'h020f008a803481d2;
        dcache[1002] = 64'h801e00ca00028040;
        dcache[1003] = 64'h827f020502c60073;
        dcache[1004] = 64'h813d02b080000057;
        dcache[1005] = 64'h005c000f0041004f;
        dcache[1006] = 64'h8007018b80928059;
        dcache[1007] = 64'h8135020402a700d1;
        dcache[1008] = 64'h012d0123813d806a;
        dcache[1009] = 64'h8088802080f80047;
        dcache[1010] = 64'h0015006200c88132;
        dcache[1011] = 64'h00e0803980408049;
        dcache[1012] = 64'h0123016181508080;
        dcache[1013] = 64'h000580ca80f40083;
        dcache[1014] = 64'h80fb805501e80007;
        dcache[1015] = 64'h013d804881468078;
        dcache[1016] = 64'h0084804580728069;
        dcache[1017] = 64'h0079010680ed010e;
        dcache[1018] = 64'h800d80dc80e1006c;
        dcache[1019] = 64'h00f380a1006a803b;
        dcache[1020] = 64'h00b100d801c4824f;
        dcache[1021] = 64'h80da8107806100b3;
        dcache[1022] = 64'h000f809b00f080a5;
        dcache[1023] = 64'h01e181c3804a0068;
        dcache[1024] = 64'h00b7014d00ca8058;
        dcache[1025] = 64'h80cc0074823400a9;
        dcache[1026] = 64'h819c00a0010200c1;
        dcache[1027] = 64'h012c825c81af00d0;
        dcache[1028] = 64'h0125010200c28042;
        dcache[1029] = 64'h00f30072816b006d;
        dcache[1030] = 64'h804a8109011780b9;
        dcache[1031] = 64'h01c481d400be8090;
        dcache[1032] = 64'h006a00d8002c0007;
        dcache[1033] = 64'h804f80ee81278017;
        dcache[1034] = 64'h8002007300c68005;
        dcache[1035] = 64'h009181b6017c8152;
        dcache[1036] = 64'h800e00f28081007b;
        dcache[1037] = 64'h8060809080df004c;
        dcache[1038] = 64'h804a006900f30027;
        dcache[1039] = 64'h8026816e006f8110;
        dcache[1040] = 64'h006400e580a1003e;
        dcache[1041] = 64'h0001808280bd0060;
        dcache[1042] = 64'h003300900048000e;
        dcache[1043] = 64'h805480be00c58103;
        dcache[1044] = 64'h0031011f80a200b0;
        dcache[1045] = 64'h805580dc807800d8;
        dcache[1046] = 64'h007700000040804c;
        dcache[1047] = 64'h800a80ae007a8089;
        dcache[1048] = 64'h0047008a801600f9;
        dcache[1049] = 64'h002c80ec802800d7;
        dcache[1050] = 64'h0089005b006580df;
        dcache[1051] = 64'h009b806800278093;
        dcache[1052] = 64'h008d011d80d900e7;
        dcache[1053] = 64'h00ba81078083005a;
        dcache[1054] = 64'h8025001e00348074;
        dcache[1055] = 64'h004000c9001980ff;
        dcache[1056] = 64'h00530155806c00be;
        dcache[1057] = 64'h801c80bc801100d4;
        dcache[1058] = 64'h001c005c0045805b;
        dcache[1059] = 64'h00b200bb80b1808b;
        dcache[1060] = 64'h805f0170000c00bb;
        dcache[1061] = 64'h814d80a600118151;
        dcache[1062] = 64'h002b00150018802a;
        dcache[1063] = 64'h00f80112812d8079;
        dcache[1064] = 64'h8026012700bd007c;
        dcache[1065] = 64'h819280850045819f;
        dcache[1066] = 64'h80740092007280fc;
        dcache[1067] = 64'h01ba004380fd8103;
        dcache[1068] = 64'h80220088011f8123;
        dcache[1069] = 64'h80ea80750052802f;
        dcache[1070] = 64'h811c0107801e80b1;
        dcache[1071] = 64'h015c0022811f8028;
        dcache[1072] = 64'h0006000c00c481cd;
        dcache[1073] = 64'h80660041801e0021;
        dcache[1074] = 64'h80a98063806b8075;
        dcache[1075] = 64'h013200008059007c;
        dcache[1076] = 64'h008c000f0054824a;
        dcache[1077] = 64'h80f98018804700b6;
        dcache[1078] = 64'h8064803f0049805b;
        dcache[1079] = 64'h015d0101002a0142;
        dcache[1080] = 64'h009f003b804081ea;
        dcache[1081] = 64'h808f804a80120058;
        dcache[1082] = 64'h8052802380228042;
        dcache[1083] = 64'h00c700fc802f00ae;
        dcache[1084] = 64'h8000007000508249;
        dcache[1085] = 64'h80b5801e8040002a;
        dcache[1086] = 64'h000280af80c18084;
        dcache[1087] = 64'h00f500c6003700d4;
        dcache[1088] = 64'h0033008580208210;
        dcache[1089] = 64'h80d9005180050013;
        dcache[1090] = 64'h0031803c80b48063;
        dcache[1091] = 64'h00c9005700b000f5;
        dcache[1092] = 64'h006300ee801881eb;
        dcache[1093] = 64'h805d0085813a8061;
        dcache[1094] = 64'h0027807b80b48051;
        dcache[1095] = 64'h001f00ed0075000d;
        dcache[1096] = 64'h0039011e8083816b;
        dcache[1097] = 64'h8056806c80bb00a3;
        dcache[1098] = 64'h80bc805100058072;
        dcache[1099] = 64'h005e003b013a0083;
        dcache[1100] = 64'h0155010b819e80a5;
        dcache[1101] = 64'h80a280eb81528043;
        dcache[1102] = 64'h00e98078801e811d;
        dcache[1103] = 64'h801d009c017b013d;
        dcache[1104] = 64'h013b014a82208091;
        dcache[1105] = 64'h803a80b480ea830c;
        dcache[1106] = 64'h00be016c00628124;
        dcache[1107] = 64'h809402c5014801ee;
        dcache[1108] = 64'h0190025d80160034;
        dcache[1109] = 64'h0146805e819f82b4;
        dcache[1110] = 64'h8080016c80380062;
        dcache[1111] = 64'h827a03120379016f;
        dcache[1112] = 64'h807e041700a50047;
        dcache[1113] = 64'h017c00f4809880f7;
        dcache[1114] = 64'h81a700b6800c814a;
        dcache[1115] = 64'h8324020d028e0066;
        dcache[1116] = 64'h80bf026480cd00f3;
        dcache[1117] = 64'h814b81550025007c;
        dcache[1118] = 64'h80e700670051808a;
        dcache[1119] = 64'h824000048071019e;
        dcache[1120] = 64'h015e00d281000010;
        dcache[1121] = 64'h8041805380af0000;
        dcache[1122] = 64'h8001006301088125;
        dcache[1123] = 64'h0164800a80b7800d;
        dcache[1124] = 64'h021f006581e88153;
        dcache[1125] = 64'h808e80aa815d004e;
        dcache[1126] = 64'h81530057027680f0;
        dcache[1127] = 64'h00f6011981468080;
        dcache[1128] = 64'h00f10057813a0086;
        dcache[1129] = 64'h80f1003c81448027;
        dcache[1130] = 64'h0097805a006d80b4;
        dcache[1131] = 64'h0195805c80b3001c;
        dcache[1132] = 64'h0069014f017a80e3;
        dcache[1133] = 64'h818d806680c080a2;
        dcache[1134] = 64'h8014805180a00027;
        dcache[1135] = 64'h0195819200040090;
        dcache[1136] = 64'h004001760059804c;
        dcache[1137] = 64'h800700638225005b;
        dcache[1138] = 64'h80bb8002009b0067;
        dcache[1139] = 64'h005b8163008080fb;
        dcache[1140] = 64'h0042012600280037;
        dcache[1141] = 64'h00cb803880888046;
        dcache[1142] = 64'h0040806400a08107;
        dcache[1143] = 64'h013d81fa007c813f;
        dcache[1144] = 64'h005a011b80340048;
        dcache[1145] = 64'h005e80d1800e8014;
        dcache[1146] = 64'h0050003901118072;
        dcache[1147] = 64'h00f681da010080af;
        dcache[1148] = 64'h00320116810f009e;
        dcache[1149] = 64'h80268081809b000d;
        dcache[1150] = 64'h8070004600e7000e;
        dcache[1151] = 64'h0018813d010880bd;
        dcache[1152] = 64'h001000bb810200ed;
        dcache[1153] = 64'h002880c480480020;
        dcache[1154] = 64'h80440026003c8067;
        dcache[1155] = 64'h807080590122810e;
        dcache[1156] = 64'h00c80171813400b4;
        dcache[1157] = 64'h005b810780008069;
        dcache[1158] = 64'h80008014007a80a0;
        dcache[1159] = 64'h004d803a00b68123;
        dcache[1160] = 64'h00660131805b008e;
        dcache[1161] = 64'h007c812e809380ff;
        dcache[1162] = 64'h0028004a00ad80a8;
        dcache[1163] = 64'h8013001600358107;
        dcache[1164] = 64'h008e0165806800df;
        dcache[1165] = 64'h00908123805381af;
        dcache[1166] = 64'h00580020007d8143;
        dcache[1167] = 64'h0031009880a880cc;
        dcache[1168] = 64'h007601fe00660089;
        dcache[1169] = 64'h80ab80a100a5834c;
        dcache[1170] = 64'h00dc802d80628079;
        dcache[1171] = 64'h807701a2809a8168;
        dcache[1172] = 64'h807802618000005a;
        dcache[1173] = 64'h8241802600398484;
        dcache[1174] = 64'h802c00ca0080806c;
        dcache[1175] = 64'h0061011c822780e5;
        dcache[1176] = 64'h806b01a200d380ab;
        dcache[1177] = 64'h818e802b000b835f;
        dcache[1178] = 64'h8003019e006b80fa;
        dcache[1179] = 64'h0176011981b68145;
        dcache[1180] = 64'h00a70071004f81ac;
        dcache[1181] = 64'h80e40060800480be;
        dcache[1182] = 64'h810c00e000308076;
        dcache[1183] = 64'h00c8014781f78159;
        dcache[1184] = 64'h0036003b005e81ba;
        dcache[1185] = 64'h8107009700418028;
        dcache[1186] = 64'h80fe0093801b8059;
        dcache[1187] = 64'h017000d18124800b;
        dcache[1188] = 64'h000b800a008e8195;
        dcache[1189] = 64'h80f4009300230055;
        dcache[1190] = 64'h801380d400108089;
        dcache[1191] = 64'h00d7004f80ac8008;
        dcache[1192] = 64'h00e0801000208264;
        dcache[1193] = 64'h8086000f80160023;
        dcache[1194] = 64'h0044802e008d0002;
        dcache[1195] = 64'h010600018027005e;
        dcache[1196] = 64'h007c0068009982fa;
        dcache[1197] = 64'h80b40067003c8066;
        dcache[1198] = 64'h801500080017005c;
        dcache[1199] = 64'h00a4009d80520062;
        dcache[1200] = 64'h009b00bf00468321;
        dcache[1201] = 64'h80e10042808e801e;
        dcache[1202] = 64'h0026003f80db8016;
        dcache[1203] = 64'h017a800a002e005d;
        dcache[1204] = 64'h00c9009c804483b2;
        dcache[1205] = 64'h8077800e81390005;
        dcache[1206] = 64'h0052007480a380ad;
        dcache[1207] = 64'h00fc000000310052;
        dcache[1208] = 64'h011100d2804d8499;
        dcache[1209] = 64'h80b3806a81a88078;
        dcache[1210] = 64'h008680a48050809d;
        dcache[1211] = 64'h017a800e0096008e;
        dcache[1212] = 64'h80e50077817283ca;
        dcache[1213] = 64'h807680f8822c80e6;
        dcache[1214] = 64'h018900c880bd8179;
        dcache[1215] = 64'h00488031012700cf;
        dcache[1216] = 64'h006b00b884748200;
        dcache[1217] = 64'h8083801d82498290;
        dcache[1218] = 64'h01250122807c8051;
        dcache[1219] = 64'h8096026301bb007e;
        dcache[1220] = 64'h01570203814b80dd;
        dcache[1221] = 64'h00a8003e80478169;
        dcache[1222] = 64'h82c8020880fa0052;
        dcache[1223] = 64'h808f01e701df001e;
        dcache[1224] = 64'h808903a8804d0280;
        dcache[1225] = 64'h808c010b81018046;
        dcache[1226] = 64'h82c001ba815b813b;
        dcache[1227] = 64'h820301d801900054;
        dcache[1228] = 64'h0021009c004200a9;
        dcache[1229] = 64'h815080a780150148;
        dcache[1230] = 64'h81490042011581c9;
        dcache[1231] = 64'h8273802e80b70063;
        dcache[1232] = 64'h019d00be81c98093;
        dcache[1233] = 64'h804b80688077000b;
        dcache[1234] = 64'h8044805701be80be;
        dcache[1235] = 64'h015000ab80e4809b;
        dcache[1236] = 64'h00dd001f81f880e9;
        dcache[1237] = 64'h817400e9806b0016;
        dcache[1238] = 64'h01038088027a81a6;
        dcache[1239] = 64'h01eb00b881e80003;
        dcache[1240] = 64'h018b0167810b803b;
        dcache[1241] = 64'h8130004d8156814c;
        dcache[1242] = 64'h000400e900c880c9;
        dcache[1243] = 64'h01338012816d8123;
        dcache[1244] = 64'h012300b3015d8176;
        dcache[1245] = 64'h816a00b381d881d4;
        dcache[1246] = 64'h8095000800ae8002;
        dcache[1247] = 64'h010a808d000580a6;
        dcache[1248] = 64'h0057027780010047;
        dcache[1249] = 64'h80a2002081fe8147;
        dcache[1250] = 64'h80fc006c008a807c;
        dcache[1251] = 64'h00c381588005811b;
        dcache[1252] = 64'h0007014e00320055;
        dcache[1253] = 64'h0168805c80d78166;
        dcache[1254] = 64'h005c000f00ab809b;
        dcache[1255] = 64'h007e814900de8225;
        dcache[1256] = 64'h003a00a7810a0071;
        dcache[1257] = 64'h0080804c803580c1;
        dcache[1258] = 64'h00120053007e8099;
        dcache[1259] = 64'h00ce80f60122806d;
        dcache[1260] = 64'h009000ec80dd8020;
        dcache[1261] = 64'h0051810680338213;
        dcache[1262] = 64'h00b0801600e780c3;
        dcache[1263] = 64'h802d805300a380a8;
        dcache[1264] = 64'h00aa800e80cf003e;
        dcache[1265] = 64'h0047811c0031825b;
        dcache[1266] = 64'h80270022006b8012;
        dcache[1267] = 64'h802f808301378059;
        dcache[1268] = 64'h014c008780c9000a;
        dcache[1269] = 64'h011e80e3804483dd;
        dcache[1270] = 64'h00478075006c8039;
        dcache[1271] = 64'h8079807200f88106;
        dcache[1272] = 64'h0144007380758010;
        dcache[1273] = 64'h00d48103805f8444;
        dcache[1274] = 64'h8030805400300001;
        dcache[1275] = 64'h805d001900478068;
        dcache[1276] = 64'h010f009900098033;
        dcache[1277] = 64'h800f812d005083fa;
        dcache[1278] = 64'h803d002200ce800c;
        dcache[1279] = 64'h0024009b0010802f;
        dcache[1280] = 64'h008301b800a4803a;
        dcache[1281] = 64'h003a003b014e8484;
        dcache[1282] = 64'h800d007a003c008b;
        dcache[1283] = 64'h806500c080218114;
        dcache[1284] = 64'h81950147003e8095;
        dcache[1285] = 64'h817700930084835e;
        dcache[1286] = 64'h808702900073007a;
        dcache[1287] = 64'h0074015e80bf80aa;
        dcache[1288] = 64'h808c00bf011a8150;
        dcache[1289] = 64'h80a100c1008f819f;
        dcache[1290] = 64'h8008026d00f10016;
        dcache[1291] = 64'h009c0161809c815f;
        dcache[1292] = 64'h00ae001400c681cc;
        dcache[1293] = 64'h804000c5008b0031;
        dcache[1294] = 64'h819b00e90006801d;
        dcache[1295] = 64'h0068013080b481d0;
        dcache[1296] = 64'h0054812400838039;
        dcache[1297] = 64'h001a8003004a002f;
        dcache[1298] = 64'h80eb008f004200b6;
        dcache[1299] = 64'h005700b800558246;
        dcache[1300] = 64'h00bf801700fa002f;
        dcache[1301] = 64'h80dd8070007a803b;
        dcache[1302] = 64'h8090001000a10156;
        dcache[1303] = 64'h0129004400a180f8;
        dcache[1304] = 64'h0068000200ea003a;
        dcache[1305] = 64'h800c807980098056;
        dcache[1306] = 64'h805e005200ed00c9;
        dcache[1307] = 64'h00ef005580108062;
        dcache[1308] = 64'h0026000901278073;
        dcache[1309] = 64'h004a009700900014;
        dcache[1310] = 64'h800d0022006c800e;
        dcache[1311] = 64'h011280010015800a;
        dcache[1312] = 64'h80818016008b8268;
        dcache[1313] = 64'h807a8054004b800c;
        dcache[1314] = 64'h805700f500d58017;
        dcache[1315] = 64'h018280a38033809b;
        dcache[1316] = 64'h802a80ad80a6823f;
        dcache[1317] = 64'h80918042806f8065;
        dcache[1318] = 64'h00a800890082808c;
        dcache[1319] = 64'h016680bd808b006a;
        dcache[1320] = 64'h000a80ab807c8499;
        dcache[1321] = 64'h801c808d81b980bb;
        dcache[1322] = 64'h004b00ee001980a4;
        dcache[1323] = 64'h012580d0000c008c;
        dcache[1324] = 64'h8138803b81c68493;
        dcache[1325] = 64'h80238054827e8011;
        dcache[1326] = 64'h0159021e80d280a4;
        dcache[1327] = 64'h802a00c8006b80ff;
        dcache[1328] = 64'h81ff80f1821f8402;
        dcache[1329] = 64'h0031809082d680cd;
        dcache[1330] = 64'h018101f382418191;
        dcache[1331] = 64'h80cd01a3024e001d;
        dcache[1332] = 64'h806f004f806981b2;
        dcache[1333] = 64'h00b300b4815b004a;
        dcache[1334] = 64'h809a00e9820580e4;
        dcache[1335] = 64'h808900d102ce80af;
        dcache[1336] = 64'h006101ee025101c3;
        dcache[1337] = 64'h00fb0076826280ca;
        dcache[1338] = 64'h813d00f181298169;
        dcache[1339] = 64'h0010030a033b004c;
        dcache[1340] = 64'h00b9812200cd016f;
        dcache[1341] = 64'h819a80c28079010c;
        dcache[1342] = 64'h8152014301930023;
        dcache[1343] = 64'h81b901ca80c781a9;
        dcache[1344] = 64'h010a007c80b580c6;
        dcache[1345] = 64'h002a005000090003;
        dcache[1346] = 64'h8014805800b4001d;
        dcache[1347] = 64'h0033009180ae8029;
        dcache[1348] = 64'h028c01f9812d813d;
        dcache[1349] = 64'h805a006f80f580b4;
        dcache[1350] = 64'h0072803802118068;
        dcache[1351] = 64'h0067809680f78007;
        dcache[1352] = 64'h01fa00aa814d8089;
        dcache[1353] = 64'h807b802c80be811d;
        dcache[1354] = 64'h00f600050165810f;
        dcache[1355] = 64'h013f805780788152;
        dcache[1356] = 64'h008a80020160802f;
        dcache[1357] = 64'h0068801981e68197;
        dcache[1358] = 64'h007a00920161812c;
        dcache[1359] = 64'h0084005200c1809e;
        dcache[1360] = 64'h0021008380230030;
        dcache[1361] = 64'h004e816a8200828a;
        dcache[1362] = 64'h80fd013001818138;
        dcache[1363] = 64'h018180a100d181ae;
        dcache[1364] = 64'h0008008d004c0059;
        dcache[1365] = 64'h00ff80d4818c8299;
        dcache[1366] = 64'h800b009e00d780d4;
        dcache[1367] = 64'h006a80bd0109818c;
        dcache[1368] = 64'h8001806d81040064;
        dcache[1369] = 64'h805780e1803d838b;
        dcache[1370] = 64'h003601160029006c;
        dcache[1371] = 64'h8002002600ed804b;
        dcache[1372] = 64'h0120805f80f08054;
        dcache[1373] = 64'h800180c8801284ba;
        dcache[1374] = 64'h00600054001b0004;
        dcache[1375] = 64'h808e004400718050;
        dcache[1376] = 64'h013080218098001a;
        dcache[1377] = 64'h00ca8062007184e8;
        dcache[1378] = 64'h8099802e00888086;
        dcache[1379] = 64'h8049808900780088;
        dcache[1380] = 64'h009980b8800b8039;
        dcache[1381] = 64'h00168049007884a0;
        dcache[1382] = 64'h8017003980068036;
        dcache[1383] = 64'h806480d5003c0064;
        dcache[1384] = 64'h010880978082001f;
        dcache[1385] = 64'h003d006000798394;
        dcache[1386] = 64'h80c08038806c015f;
        dcache[1387] = 64'h805c806e00b300cc;
        dcache[1388] = 64'h017580df00300013;
        dcache[1389] = 64'h003600bc01458231;
        dcache[1390] = 64'h80a98091805c0146;
        dcache[1391] = 64'h0026003900f7004a;
        dcache[1392] = 64'h0036801700af0017;
        dcache[1393] = 64'h8044024e01b98144;
        dcache[1394] = 64'h807480cb80ca012b;
        dcache[1395] = 64'h80350139003b0004;
        dcache[1396] = 64'h817c805f00d780e9;
        dcache[1397] = 64'h80b30254014f80fc;
        dcache[1398] = 64'h802100a1811d00b0;
        dcache[1399] = 64'h80b5015900d9805b;
        dcache[1400] = 64'h811c805d0158810e;
        dcache[1401] = 64'h80f600dd014b8062;
        dcache[1402] = 64'h80d9020c005b004c;
        dcache[1403] = 64'h800a019700a480e8;
        dcache[1404] = 64'h00d48013012780df;
        dcache[1405] = 64'h804c809c00430080;
        dcache[1406] = 64'h8155011a00ab00d2;
        dcache[1407] = 64'h802a01000070817c;
        dcache[1408] = 64'h00d5807500bd8031;
        dcache[1409] = 64'h002d806c0040007a;
        dcache[1410] = 64'h80b2001600fa00fe;
        dcache[1411] = 64'h0025004580328174;
        dcache[1412] = 64'h0082001a014300ae;
        dcache[1413] = 64'h802680c400278060;
        dcache[1414] = 64'h80410030014400bc;
        dcache[1415] = 64'h0081001480158109;
        dcache[1416] = 64'h0005002301040106;
        dcache[1417] = 64'h8059805300b2805e;
        dcache[1418] = 64'h80a2803b01b20076;
        dcache[1419] = 64'h011a000f8050808f;
        dcache[1420] = 64'h8052806f01988004;
        dcache[1421] = 64'h00c5800600d48085;
        dcache[1422] = 64'h0046800500590011;
        dcache[1423] = 64'h01a8801000518027;
        dcache[1424] = 64'h806c800480248069;
        dcache[1425] = 64'h007d8041801980d3;
        dcache[1426] = 64'h009c00730055003c;
        dcache[1427] = 64'h012a805100d88044;
        dcache[1428] = 64'h002280de80db80d9;
        dcache[1429] = 64'h00f3802980b28033;
        dcache[1430] = 64'h01af003400960009;
        dcache[1431] = 64'h002380d600988096;
        dcache[1432] = 64'h000580fa829781b0;
        dcache[1433] = 64'h804080518092804b;
        dcache[1434] = 64'h016d00ad00ea8015;
        dcache[1435] = 64'h0052813c806c80a2;
        dcache[1436] = 64'h81f0824482418229;
        dcache[1437] = 64'h80aa81278252804d;
        dcache[1438] = 64'h01df01bb00220059;
        dcache[1439] = 64'h803700ed00de8107;
        dcache[1440] = 64'h81b782ad806b82f9;
        dcache[1441] = 64'h006f00f18206004f;
        dcache[1442] = 64'h0423803181a68107;
        dcache[1443] = 64'h80d6804780ad8008;
        dcache[1444] = 64'h808100320057821c;
        dcache[1445] = 64'h00ec01b780bb01ea;
        dcache[1446] = 64'h8097803e82df824e;
        dcache[1447] = 64'h00508053008b80c4;
        dcache[1448] = 64'h0194005d005200b9;
        dcache[1449] = 64'h0273000b807900d4;
        dcache[1450] = 64'h81f380a081fb81c8;
        dcache[1451] = 64'h0081019801fb80b3;
        dcache[1452] = 64'h0038806e803a013a;
        dcache[1453] = 64'h80dd803d001380c7;
        dcache[1454] = 64'h81b000c101d58175;
        dcache[1455] = 64'h81448091815580f1;
        dcache[1456] = 64'h000b800800ce00ea;
        dcache[1457] = 64'h80c500fe802d00e1;
        dcache[1458] = 64'h003200ef006180be;
        dcache[1459] = 64'h813e00c7814c8075;
        dcache[1460] = 64'h019100c780778098;
        dcache[1461] = 64'h001c0007804880fb;
        dcache[1462] = 64'h00ea006501800014;
        dcache[1463] = 64'h80800099006c804e;
        dcache[1464] = 64'h01ce00d9813c816a;
        dcache[1465] = 64'h8081807580d780d0;
        dcache[1466] = 64'h00f000cf01598184;
        dcache[1467] = 64'h00de80cb8115810f;
        dcache[1468] = 64'h8079802c016e009b;
        dcache[1469] = 64'h0059802080d88251;
        dcache[1470] = 64'h00bb01390176817b;
        dcache[1471] = 64'h008f006100938014;
        dcache[1472] = 64'h002781bb81360010;
        dcache[1473] = 64'h8049817f80d28400;
        dcache[1474] = 64'h8026018000fe801d;
        dcache[1475] = 64'h01ce80140090812b;
        dcache[1476] = 64'h00368092816a8054;
        dcache[1477] = 64'h00618026816e8491;
        dcache[1478] = 64'h805d007100520005;
        dcache[1479] = 64'h800b80840019801d;
        dcache[1480] = 64'h00ef8123816d803f;
        dcache[1481] = 64'h806f8003007c841b;
        dcache[1482] = 64'h00140034002b000e;
        dcache[1483] = 64'h8053804480d0005d;
        dcache[1484] = 64'h0183814680db801d;
        dcache[1485] = 64'h80168032011f8387;
        dcache[1486] = 64'h8041002f80c7803c;
        dcache[1487] = 64'h8002006a007d0062;
        dcache[1488] = 64'h007d80ec003b809c;
        dcache[1489] = 64'h002a009800778234;
        dcache[1490] = 64'h803f80b780770024;
        dcache[1491] = 64'h0010800d00b30098;
        dcache[1492] = 64'h009d80d6001e80b5;
        dcache[1493] = 64'h005400b4002781ee;
        dcache[1494] = 64'h809e80f080a00063;
        dcache[1495] = 64'h000e002100ac008d;
        dcache[1496] = 64'h018780f08107805b;
        dcache[1497] = 64'h002e00e500d88073;
        dcache[1498] = 64'h808580bf80b100a2;
        dcache[1499] = 64'h00138068015a00aa;
        dcache[1500] = 64'h015f81478051803e;
        dcache[1501] = 64'h005c0134014e0029;
        dcache[1502] = 64'h8045811f80a30057;
        dcache[1503] = 64'h801300dc01ea0075;
        dcache[1504] = 64'h803a8172006e80a1;
        dcache[1505] = 64'h80450283016c002f;
        dcache[1506] = 64'h0018809981820095;
        dcache[1507] = 64'h810c0177022e8017;
        dcache[1508] = 64'h825880ed01438120;
        dcache[1509] = 64'h801d010e01080079;
        dcache[1510] = 64'h805c014980af003c;
        dcache[1511] = 64'h80ac00f101dd8036;
        dcache[1512] = 64'h8081800601ed8061;
        dcache[1513] = 64'h80480054008c0056;
        dcache[1514] = 64'h805b019d80510020;
        dcache[1515] = 64'h8005013400bb0007;
        dcache[1516] = 64'h00128063014b805c;
        dcache[1517] = 64'h0046001200ab0078;
        dcache[1518] = 64'h801000c9010700c3;
        dcache[1519] = 64'h80f1013700e68079;
        dcache[1520] = 64'h007200860150806e;
        dcache[1521] = 64'h0067808800e40004;
        dcache[1522] = 64'h80ef005501810149;
        dcache[1523] = 64'h80810031006a8109;
        dcache[1524] = 64'h002100a1018f007d;
        dcache[1525] = 64'h80018027008c8047;
        dcache[1526] = 64'h8083800b010400fb;
        dcache[1527] = 64'h80068045001c80f1;
        dcache[1528] = 64'h001d00b600e40015;
        dcache[1529] = 64'h0027003f00bc8077;
        dcache[1530] = 64'h801e8037012f00ba;
        dcache[1531] = 64'h0080804d00bf8092;
        dcache[1532] = 64'h80cb80ed8039001e;
        dcache[1533] = 64'h00bc802c00528061;
        dcache[1534] = 64'h0070803c007d00cf;
        dcache[1535] = 64'h00a1800a015e8054;
        dcache[1536] = 64'h0090807e805a0032;
        dcache[1537] = 64'h017b806b80470031;
        dcache[1538] = 64'h008d800900420015;
        dcache[1539] = 64'h00a5002100f48045;
        dcache[1540] = 64'h008c80c9822a000c;
        dcache[1541] = 64'h00ee803f80108003;
        dcache[1542] = 64'h00c4001400a4002f;
        dcache[1543] = 64'h00ab803a8012807b;
        dcache[1544] = 64'h8006810f82ae003b;
        dcache[1545] = 64'h004c806d81208029;
        dcache[1546] = 64'h01e080350090801c;
        dcache[1547] = 64'h001b8088004e8143;
        dcache[1548] = 64'h813381ff8244000a;
        dcache[1549] = 64'h80ec00c1810c00d3;
        dcache[1550] = 64'h020e011400bc0014;
        dcache[1551] = 64'h80b78035806380ff;
        dcache[1552] = 64'h80a98123807b000b;
        dcache[1553] = 64'h801c0152802800d6;
        dcache[1554] = 64'h01eb001880b28111;
        dcache[1555] = 64'h802f80e881118006;
        dcache[1556] = 64'h005d80a5011780f4;
        dcache[1557] = 64'h00ab012980680201;
        dcache[1558] = 64'h00d6812981f48240;
        dcache[1559] = 64'h800c80cf802f0009;
        dcache[1560] = 64'h00ce021201b3806d;
        dcache[1561] = 64'h02fb014600fa0127;
        dcache[1562] = 64'h811e82a6821b835f;
        dcache[1563] = 64'h801e810d00c90018;
        dcache[1564] = 64'h806a00d2016a005e;
        dcache[1565] = 64'h01a6017001820091;
        dcache[1566] = 64'h008f817a0089812b;
        dcache[1567] = 64'h8058820780f80073;
        dcache[1568] = 64'h00b80118811b012b;
        dcache[1569] = 64'h00c000ae80288032;
        dcache[1570] = 64'h00d1001780bd8138;
        dcache[1571] = 64'h80e601070071007a;
        dcache[1572] = 64'h00f901ae0004812e;
        dcache[1573] = 64'h803d805080778100;
        dcache[1574] = 64'h808000a500a300bd;
        dcache[1575] = 64'h806b806e002580a2;
        dcache[1576] = 64'h020d025c8160817e;
        dcache[1577] = 64'h810d002180c180cc;
        dcache[1578] = 64'h8020004b020480fa;
        dcache[1579] = 64'h00ed00918169002c;
        dcache[1580] = 64'h805980bb018e002e;
        dcache[1581] = 64'h01590128002f8213;
        dcache[1582] = 64'h0098016300d38138;
        dcache[1583] = 64'h0114000500910033;
        dcache[1584] = 64'h00b9817980d080b0;
        dcache[1585] = 64'h00f8806300688223;
        dcache[1586] = 64'h8036006680f50099;
        dcache[1587] = 64'h00bf808e8032000f;
        dcache[1588] = 64'h015d83918151826d;
        dcache[1589] = 64'h008e008e80de8235;
        dcache[1590] = 64'h801f801e802c00aa;
        dcache[1591] = 64'h00188063806f00d5;
        dcache[1592] = 64'h00f8837380628125;
        dcache[1593] = 64'h009b00a38012811a;
        dcache[1594] = 64'h000200158041002f;
        dcache[1595] = 64'h800f8120001b0083;
        dcache[1596] = 64'h00fc829c80578023;
        dcache[1597] = 64'h00ac004401178012;
        dcache[1598] = 64'h8014808b815d806a;
        dcache[1599] = 64'h00ae803f00670081;
        dcache[1600] = 64'h00f7823e80358019;
        dcache[1601] = 64'h802a00c600d20031;
        dcache[1602] = 64'h804580bb81210045;
        dcache[1603] = 64'h004b001d00698015;
        dcache[1604] = 64'h00fd8211808c804d;
        dcache[1605] = 64'h001000d600980092;
        dcache[1606] = 64'h80318072814700a6;
        dcache[1607] = 64'h8043004780180000;
        dcache[1608] = 64'h00e280eb811b8016;
        dcache[1609] = 64'h80240060009800e6;
        dcache[1610] = 64'h0048800a808e8027;
        dcache[1611] = 64'h8073002e0111809b;
        dcache[1612] = 64'h006981958066809d;
        dcache[1613] = 64'h002f00d9011a00c4;
        dcache[1614] = 64'h00ec80aa8066002e;
        dcache[1615] = 64'h80cb005501c88055;
        dcache[1616] = 64'h8177819a002a80a4;
        dcache[1617] = 64'h80ce01c901190079;
        dcache[1618] = 64'h0043805580c1008d;
        dcache[1619] = 64'h807b009301c08051;
        dcache[1620] = 64'h819080f501a78131;
        dcache[1621] = 64'h0016011e00b70097;
        dcache[1622] = 64'h004e007580198052;
        dcache[1623] = 64'h805000c30163001b;
        dcache[1624] = 64'h8042801b019c8046;
        dcache[1625] = 64'h003600e3006700b3;
        dcache[1626] = 64'h802b00a200018012;
        dcache[1627] = 64'h80d2013900dd005c;
        dcache[1628] = 64'h80118019014e805a;
        dcache[1629] = 64'h00aa003d00b30065;
        dcache[1630] = 64'h80800068008e0120;
        dcache[1631] = 64'h808e005d0087003d;
        dcache[1632] = 64'h0064001701328032;
        dcache[1633] = 64'h00e8003a01620044;
        dcache[1634] = 64'h80a4005c012001a3;
        dcache[1635] = 64'h80aa80430053810a;
        dcache[1636] = 64'h01060034011480ea;
        dcache[1637] = 64'h0052801401390057;
        dcache[1638] = 64'h8065804e00b10120;
        dcache[1639] = 64'h0074009300ab8113;
        dcache[1640] = 64'h0044005f80118024;
        dcache[1641] = 64'h0099006000d08019;
        dcache[1642] = 64'h80048000016400a1;
        dcache[1643] = 64'h01248011010080a0;
        dcache[1644] = 64'h00e4800a80fc8037;
        dcache[1645] = 64'h013f001700df0022;
        dcache[1646] = 64'h0096805b007300d5;
        dcache[1647] = 64'h010b802d801c8102;
        dcache[1648] = 64'h0082807481900062;
        dcache[1649] = 64'h00b08067002d00c0;
        dcache[1650] = 64'h0085006080f50074;
        dcache[1651] = 64'h011480618079806f;
        dcache[1652] = 64'h8036801981ff800c;
        dcache[1653] = 64'h002480a980bd00df;
        dcache[1654] = 64'h00e2008280eb00d6;
        dcache[1655] = 64'h00c080858044802b;
        dcache[1656] = 64'h00f080af81b000f4;
        dcache[1657] = 64'h0005007f808b0044;
        dcache[1658] = 64'h0093801c003600a3;
        dcache[1659] = 64'h8063811b8084816f;
        dcache[1660] = 64'h00c9800781ad0085;
        dcache[1661] = 64'h818600a58006003e;
        dcache[1662] = 64'h0081005c01748041;
        dcache[1663] = 64'h0055001b815e807a;
        dcache[1664] = 64'h8002000b80c100e4;
        dcache[1665] = 64'h81360118008d007a;
        dcache[1666] = 64'h008f0097008c8090;
        dcache[1667] = 64'h002700e8814b0005;
        dcache[1668] = 64'h001f803f016f0007;
        dcache[1669] = 64'h001b017d023800c9;
        dcache[1670] = 64'h01cf80f9801480f6;
        dcache[1671] = 64'h80b5819080ab80e2;
        dcache[1672] = 64'h814f010702bd8119;
        dcache[1673] = 64'h033002b702bc0119;
        dcache[1674] = 64'h811282d6803d8393;
        dcache[1675] = 64'h012b8282001800f4;
        dcache[1676] = 64'h8084003000a00026;
        dcache[1677] = 64'h01b301c401660129;
        dcache[1678] = 64'h80168179800a815f;
        dcache[1679] = 64'h0113814f815b00dc;
        dcache[1680] = 64'h00da0096813800da;
        dcache[1681] = 64'h007f008780900044;
        dcache[1682] = 64'h0081004d80c28155;
        dcache[1683] = 64'h80c700bf00dd0059;
        dcache[1684] = 64'h004900ee005080ea;
        dcache[1685] = 64'h8139802f0042801b;
        dcache[1686] = 64'h80d400e5004a00be;
        dcache[1687] = 64'h0094004100f580c9;
        dcache[1688] = 64'h029d01e60074813d;
        dcache[1689] = 64'h806f02b4815f80ae;
        dcache[1690] = 64'h00648212004c020f;
        dcache[1691] = 64'h820c01d880f6822b;
        dcache[1692] = 64'h006d810f0156804d;
        dcache[1693] = 64'h01ab014e011b80df;
        dcache[1694] = 64'h00c580ac80e180b8;
        dcache[1695] = 64'h0030001c00928103;
        dcache[1696] = 64'h00ee820a80d68146;
        dcache[1697] = 64'h007d00a100c38003;
        dcache[1698] = 64'h80cd80a981a3802b;
        dcache[1699] = 64'h018480b580270052;
        dcache[1700] = 64'h002384258096816f;
        dcache[1701] = 64'h007c006c00a3006c;
        dcache[1702] = 64'h0038801181900083;
        dcache[1703] = 64'h0123810580760156;
        dcache[1704] = 64'h0149836f000880b9;
        dcache[1705] = 64'h0124009000980151;
        dcache[1706] = 64'h801900728137007e;
        dcache[1707] = 64'h005780bb809f00bc;
        dcache[1708] = 64'h0085830d80388090;
        dcache[1709] = 64'h00150046001b00ca;
        dcache[1710] = 64'h00ec800280e5006e;
        dcache[1711] = 64'h0057802180c2002c;
        dcache[1712] = 64'h00e68266000a8020;
        dcache[1713] = 64'h004b002d005100e1;
        dcache[1714] = 64'h00d4804e81b8001e;
        dcache[1715] = 64'h8094006600308010;
        dcache[1716] = 64'h00b38191801b001b;
        dcache[1717] = 64'h00700051009400b3;
        dcache[1718] = 64'h0153803e8199806b;
        dcache[1719] = 64'h80ae00970061804d;
        dcache[1720] = 64'h00d8816d8103802c;
        dcache[1721] = 64'h00228036010e00d8;
        dcache[1722] = 64'h013d809a80ea0060;
        dcache[1723] = 64'h8054004200878081;
        dcache[1724] = 64'h801a810a80628023;
        dcache[1725] = 64'h80b1007c00df00c9;
        dcache[1726] = 64'h014d8036804a0097;
        dcache[1727] = 64'h80fa001501768087;
        dcache[1728] = 64'h815380a5001b802f;
        dcache[1729] = 64'h8045011000ec008b;
        dcache[1730] = 64'h00d40070806d0078;
        dcache[1731] = 64'h816d005b014c8061;
        dcache[1732] = 64'h816880c601538092;
        dcache[1733] = 64'h007b015e003900a7;
        dcache[1734] = 64'h000a00e200948028;
        dcache[1735] = 64'h80ec001a00c38059;
        dcache[1736] = 64'h8091807201f48063;
        dcache[1737] = 64'h005101910020006f;
        dcache[1738] = 64'h806f000d010b0083;
        dcache[1739] = 64'h80f60032009b8086;
        dcache[1740] = 64'h00290072013e000a;
        dcache[1741] = 64'h00fc007901600085;
        dcache[1742] = 64'h80dd003b017300fa;
        dcache[1743] = 64'h8013801a011a0018;
        dcache[1744] = 64'h003f805e0181004c;
        dcache[1745] = 64'h010300ed01ef0035;
        dcache[1746] = 64'h8127000300c70124;
        dcache[1747] = 64'h808c801200bc8079;
        dcache[1748] = 64'h012c0020804a8037;
        dcache[1749] = 64'h00530011015e805c;
        dcache[1750] = 64'h0026804201230161;
        dcache[1751] = 64'h00a7000700eb80f3;
        dcache[1752] = 64'h00e3007b81a78013;
        dcache[1753] = 64'h00a2003700b50040;
        dcache[1754] = 64'h00850060007d002e;
        dcache[1755] = 64'h0154007d006e80c3;
        dcache[1756] = 64'h009f008a81a8807c;
        dcache[1757] = 64'h009c0037007c0056;
        dcache[1758] = 64'h0072000b80320082;
        dcache[1759] = 64'h012280d680908133;
        dcache[1760] = 64'h00ab00ca81320020;
        dcache[1761] = 64'h800680a280158088;
        dcache[1762] = 64'h003800cf80e800fd;
        dcache[1763] = 64'h01f8814b811a8081;
        dcache[1764] = 64'h0054004a80ff0000;
        dcache[1765] = 64'h806d006f80e20099;
        dcache[1766] = 64'h005300c280fd008a;
        dcache[1767] = 64'h00a9812280fa807a;
        dcache[1768] = 64'h01960056004280b6;
        dcache[1769] = 64'h80b2803f8070001c;
        dcache[1770] = 64'h003b803c801b019e;
        dcache[1771] = 64'h0109808980ad80cc;
        dcache[1772] = 64'h0103804980680065;
        dcache[1773] = 64'h818300b0010d0040;
        dcache[1774] = 64'h802a0065802a0133;
        dcache[1775] = 64'h00720031805b8010;
        dcache[1776] = 64'h80f100d8007a011f;
        dcache[1777] = 64'h81160128013400f1;
        dcache[1778] = 64'h005300c100768054;
        dcache[1779] = 64'h00a58000807f00b4;
        dcache[1780] = 64'h811f8028012801c9;
        dcache[1781] = 64'h008b0200019e8025;
        dcache[1782] = 64'h0327801e0113804f;
        dcache[1783] = 64'h81a681178059812f;
        dcache[1784] = 64'h00580124022b80d5;
        dcache[1785] = 64'h0376015c010d0097;
        dcache[1786] = 64'h8108830381d88131;
        dcache[1787] = 64'h00ec818700de01cf;
        dcache[1788] = 64'h00740133021e0051;
        dcache[1789] = 64'h01fc01f101c200da;
        dcache[1790] = 64'h80d9824000af81c2;
        dcache[1791] = 64'h0183819080a70135;
        dcache[1792] = 64'h0083002b002f80c5;
        dcache[1793] = 64'h80058042800d8044;
        dcache[1794] = 64'h808580ad00d280a2;
        dcache[1795] = 64'h00ae80918077001c;
        dcache[1796] = 64'h000b012b013580c6;
        dcache[1797] = 64'h81b700c480d58041;
        dcache[1798] = 64'h81b80194804b0103;
        dcache[1799] = 64'h00f780b3016f80fa;
        dcache[1800] = 64'h01850251016281ec;
        dcache[1801] = 64'h80830104803e01be;
        dcache[1802] = 64'h8075808e00d200da;
        dcache[1803] = 64'h000180f1805d8026;
        dcache[1804] = 64'h003a807000ce004a;
        dcache[1805] = 64'h00e902460076015c;
        dcache[1806] = 64'h002680ce816180a1;
        dcache[1807] = 64'h00620058005e005a;
        dcache[1808] = 64'h80cf81e0801e813f;
        dcache[1809] = 64'h80ba010800d500d2;
        dcache[1810] = 64'h80bc8019811900a0;
        dcache[1811] = 64'h02a880ad8017004c;
        dcache[1812] = 64'h8006820880d80020;
        dcache[1813] = 64'h004000a801440135;
        dcache[1814] = 64'h003300e1814000b3;
        dcache[1815] = 64'h00cc807681380034;
        dcache[1816] = 64'h00c281f080018110;
        dcache[1817] = 64'h00f2009f00480178;
        dcache[1818] = 64'h0050005080b20051;
        dcache[1819] = 64'h0059004d8145803a;
        dcache[1820] = 64'h014081dc00168113;
        dcache[1821] = 64'h003b002c009000f0;
        dcache[1822] = 64'h010a00968198004a;
        dcache[1823] = 64'h006b811c81528031;
        dcache[1824] = 64'h013b82050046810c;
        dcache[1825] = 64'h00c4802500c40043;
        dcache[1826] = 64'h0201009e828b006d;
        dcache[1827] = 64'h8035804c805e804d;
        dcache[1828] = 64'h0119814b00c38062;
        dcache[1829] = 64'h803d003c001e0090;
        dcache[1830] = 64'h01ea003c815a000d;
        dcache[1831] = 64'h80af80ce801d0054;
        dcache[1832] = 64'h001680c6800b8004;
        dcache[1833] = 64'h8013800700a200cc;
        dcache[1834] = 64'h01640043807f8044;
        dcache[1835] = 64'h805f80c60060002d;
        dcache[1836] = 64'h80c180bb80a30032;
        dcache[1837] = 64'h805b00cf00e20062;
        dcache[1838] = 64'h01ae00d300d0007c;
        dcache[1839] = 64'h810980d000790002;
        dcache[1840] = 64'h80f0000c00528093;
        dcache[1841] = 64'h00cb0084007d0089;
        dcache[1842] = 64'h00f3802300570016;
        dcache[1843] = 64'h80f88046011e001e;
        dcache[1844] = 64'h816800b901498067;
        dcache[1845] = 64'h0109013900430153;
        dcache[1846] = 64'h809d004c0061003e;
        dcache[1847] = 64'h80c88012010c001f;
        dcache[1848] = 64'h8013804f0122005a;
        dcache[1849] = 64'h006b0185008b00a3;
        dcache[1850] = 64'h807f803e019900b0;
        dcache[1851] = 64'h80c1800900c98077;
        dcache[1852] = 64'h00cc006500408086;
        dcache[1853] = 64'h013b013601468004;
        dcache[1854] = 64'h80358097009e00a6;
        dcache[1855] = 64'h80390016010d804d;
        dcache[1856] = 64'h00c8000e009e8072;
        dcache[1857] = 64'h012c009a01c7803a;
        dcache[1858] = 64'h006d002e012f0051;
        dcache[1859] = 64'h800a001600878052;
        dcache[1860] = 64'h018300b1810080a0;
        dcache[1861] = 64'h00fa0067016f0009;
        dcache[1862] = 64'h009f802800220048;
        dcache[1863] = 64'h01a8800e00e6804a;
        dcache[1864] = 64'h0086008080c9805f;
        dcache[1865] = 64'h0089009b00e48028;
        dcache[1866] = 64'h00940050803e0109;
        dcache[1867] = 64'h01aa80c9802a80ce;
        dcache[1868] = 64'h0096016b80b58007;
        dcache[1869] = 64'h0076010d00010066;
        dcache[1870] = 64'h008a003b810300e7;
        dcache[1871] = 64'h019b80fd811480de;
        dcache[1872] = 64'h00d10087807c0042;
        dcache[1873] = 64'h8032007e807b805a;
        dcache[1874] = 64'h00b2000a80980136;
        dcache[1875] = 64'h016f805f80ef8129;
        dcache[1876] = 64'h012e00d6002b0059;
        dcache[1877] = 64'h800100cb00600001;
        dcache[1878] = 64'h00c480ab80970040;
        dcache[1879] = 64'h005180f4813f8090;
        dcache[1880] = 64'h00c9008800870077;
        dcache[1881] = 64'h801a009000f68040;
        dcache[1882] = 64'h00988016811400a3;
        dcache[1883] = 64'h00b180fd805f8130;
        dcache[1884] = 64'h0015008a00c800f7;
        dcache[1885] = 64'h80de015400dd801a;
        dcache[1886] = 64'h0043803980f4003d;
        dcache[1887] = 64'h002480fc804080de;
        dcache[1888] = 64'h80cf00700180013d;
        dcache[1889] = 64'h80ee024900f7002b;
        dcache[1890] = 64'h806200e18015009d;
        dcache[1891] = 64'h005081018074804f;
        dcache[1892] = 64'h8199005501bf036a;
        dcache[1893] = 64'h01fc035401c880a7;
        dcache[1894] = 64'h03eb802f000280e3;
        dcache[1895] = 64'h8085823e80b9810c;
        dcache[1896] = 64'h820700b902ae01a3;
        dcache[1897] = 64'h0238028502630047;
        dcache[1898] = 64'h810281c380ff8267;
        dcache[1899] = 64'h0152821280940002;
        dcache[1900] = 64'h80ad015902198018;
        dcache[1901] = 64'h017d01c801f400da;
        dcache[1902] = 64'h80b781d400bb81ee;
        dcache[1903] = 64'h024180c880bd0136;
        dcache[1904] = 64'h801e802a803d804b;
        dcache[1905] = 64'h0011804d0031803d;
        dcache[1906] = 64'h80058023001b0052;
        dcache[1907] = 64'h003c00290003003b;
        dcache[1908] = 64'h003e00e5014c80d8;
        dcache[1909] = 64'h81510117808800a3;
        dcache[1910] = 64'h81180134805e0109;
        dcache[1911] = 64'h0043002b0091817c;
        dcache[1912] = 64'h01b601ee018b8255;
        dcache[1913] = 64'h012a019680090239;
        dcache[1914] = 64'h00d7819d00cf008f;
        dcache[1915] = 64'h80c180e6000280c3;
        dcache[1916] = 64'h8047004000190167;
        dcache[1917] = 64'h00a40162000100d2;
        dcache[1918] = 64'h804f8017808500de;
        dcache[1919] = 64'h003f802c01bd00db;
        dcache[1920] = 64'h00cc800d801f8005;
        dcache[1921] = 64'h805200d0800c00b1;
        dcache[1922] = 64'h805d810281f70076;
        dcache[1923] = 64'h018901140083804f;
        dcache[1924] = 64'h00b18000804c0028;
        dcache[1925] = 64'h803000d600ed00bc;
        dcache[1926] = 64'h80030036817a0015;
        dcache[1927] = 64'h00ec00a880fc801a;
        dcache[1928] = 64'h00838022802c8081;
        dcache[1929] = 64'h00f10027002b00fe;
        dcache[1930] = 64'h007d00d9826b80a2;
        dcache[1931] = 64'h0030000780488037;
        dcache[1932] = 64'h00cb8049000780c2;
        dcache[1933] = 64'h0032005f8003007c;
        dcache[1934] = 64'h010c007c83c4007f;
        dcache[1935] = 64'h007180a1807d8079;
        dcache[1936] = 64'h0022809600398038;
        dcache[1937] = 64'h0068803200aa004f;
        dcache[1938] = 64'h01d500ca82a80017;
        dcache[1939] = 64'h806280b5811f8068;
        dcache[1940] = 64'h008980f9004c8078;
        dcache[1941] = 64'h80188049803a0080;
        dcache[1942] = 64'h025c002180d8802c;
        dcache[1943] = 64'h8074806b807e8004;
        dcache[1944] = 64'h0066807f804f8049;
        dcache[1945] = 64'h801b803100a70025;
        dcache[1946] = 64'h0208007b00e98041;
        dcache[1947] = 64'h80c580a58087002d;
        dcache[1948] = 64'h815c002980738016;
        dcache[1949] = 64'h0074005d00730043;
        dcache[1950] = 64'h015e007901018012;
        dcache[1951] = 64'h80e90009000a0033;
        dcache[1952] = 64'h818e800e003480ba;
        dcache[1953] = 64'h01580047002300ae;
        dcache[1954] = 64'h0061002900d88051;
        dcache[1955] = 64'h805d0013003e002f;
        dcache[1956] = 64'h80df801400d580fd;
        dcache[1957] = 64'h014200a700a500b3;
        dcache[1958] = 64'h8061800001018030;
        dcache[1959] = 64'h80d50034002080ac;
        dcache[1960] = 64'h00b28066006b8012;
        dcache[1961] = 64'h00e200e500d1009c;
        dcache[1962] = 64'h8078802201410014;
        dcache[1963] = 64'h80af00fd001b80a7;
        dcache[1964] = 64'h018f803b80328032;
        dcache[1965] = 64'h00a1009502000035;
        dcache[1966] = 64'h8014000700f40061;
        dcache[1967] = 64'h8046003f00e28001;
        dcache[1968] = 64'h00db8021002f80c0;
        dcache[1969] = 64'h007b00f701688039;
        dcache[1970] = 64'h008d801400b500c7;
        dcache[1971] = 64'h006c005c0101803e;
        dcache[1972] = 64'h00b1001180df804f;
        dcache[1973] = 64'h007700eb00bf803a;
        dcache[1974] = 64'h0053006d002700e3;
        dcache[1975] = 64'h01a9804700648044;
        dcache[1976] = 64'h00ba800a80d5007f;
        dcache[1977] = 64'h00ad01730054002e;
        dcache[1978] = 64'h00230080802200e2;
        dcache[1979] = 64'h00ea803b8089813f;
        dcache[1980] = 64'h806e006e803f0039;
        dcache[1981] = 64'h001700a380de0020;
        dcache[1982] = 64'h001000b5804000b1;
        dcache[1983] = 64'h00d9808480c4807d;
        dcache[1984] = 64'h004a001f80610067;
        dcache[1985] = 64'h0016007b80ad8097;
        dcache[1986] = 64'h00af804580860076;
        dcache[1987] = 64'h00b700048025809f;
        dcache[1988] = 64'h004a0059002300eb;
        dcache[1989] = 64'h800c00e700ff809b;
        dcache[1990] = 64'h002c80b78019006d;
        dcache[1991] = 64'h00608037801e80cb;
        dcache[1992] = 64'h00860031003f00d5;
        dcache[1993] = 64'h80a8009b800a80d5;
        dcache[1994] = 64'h0043804c80230009;
        dcache[1995] = 64'h00b180c681148048;
        dcache[1996] = 64'h80780046006a006f;
        dcache[1997] = 64'h811c01088059812b;
        dcache[1998] = 64'h804b803080fd0086;
        dcache[1999] = 64'h80308011800480bb;
        dcache[2000] = 64'h80ab806600c2002c;
        dcache[2001] = 64'h80708069808c804e;
        dcache[2002] = 64'h00b100cb00a58061;
        dcache[2003] = 64'h8064000e801d80fe;
        dcache[2004] = 64'h814a015900a1024c;
        dcache[2005] = 64'h022200f30159805c;
        dcache[2006] = 64'h020080ff013f8197;
        dcache[2007] = 64'h0111813180fc8003;
        dcache[2008] = 64'h819b00b2016700f1;
        dcache[2009] = 64'h00df0010002c0077;
        dcache[2010] = 64'h814880e6017a81ca;
        dcache[2011] = 64'h01b1804c812280b9;
        dcache[2012] = 64'h8137019c020b807a;
        dcache[2013] = 64'h808280e3017c017c;
        dcache[2014] = 64'h00e7800e007681c5;
        dcache[2015] = 64'h014281308066012f;
        dcache[2016] = 64'h010e00b2810f8019;
        dcache[2017] = 64'h80b6817981170032;
        dcache[2018] = 64'h80970109012b8137;
        dcache[2019] = 64'h014a817280b20062;
        dcache[2020] = 64'h802c00a4010c0076;
        dcache[2021] = 64'h81090160808b8001;
        dcache[2022] = 64'h80c400c60001013f;
        dcache[2023] = 64'h006980ab81070013;
        dcache[2024] = 64'h022c027d009e811f;
        dcache[2025] = 64'h001b001080550109;
        dcache[2026] = 64'h801a802901970098;
        dcache[2027] = 64'h80b00003001080dd;
        dcache[2028] = 64'h003d025c00ac0083;
        dcache[2029] = 64'h002400f50122020c;
        dcache[2030] = 64'h81d7808a80f201df;
        dcache[2031] = 64'h008580d900908095;
        dcache[2032] = 64'h8004012a001700e7;
        dcache[2033] = 64'h004701220197000f;
        dcache[2034] = 64'h0081818982af0038;
        dcache[2035] = 64'h008300ed00ad0003;
        dcache[2036] = 64'h00380166002f001f;
        dcache[2037] = 64'h0042012a00af00ba;
        dcache[2038] = 64'h004b80db82468062;
        dcache[2039] = 64'h0116805e800e808e;
        dcache[2040] = 64'h8046010c00220023;
        dcache[2041] = 64'h01000024807e0053;
        dcache[2042] = 64'h00ad80398379801c;
        dcache[2043] = 64'h00a00034007080ad;
        dcache[2044] = 64'h805b006580108043;
        dcache[2045] = 64'h00c00055805a0083;
        dcache[2046] = 64'h0167009282ef8070;
        dcache[2047] = 64'h003f806380b68007;
        dcache[2048] = 64'h80e60113802580fc;
        dcache[2049] = 64'h8008001180890038;
        dcache[2050] = 64'h01a3003082178041;
        dcache[2051] = 64'h802d8076814e802f;
        dcache[2052] = 64'h80eb001b801a81cf;
        dcache[2053] = 64'h8061800a805a0018;
        dcache[2054] = 64'h0226001c00548008;
        dcache[2055] = 64'h806680aa8165808b;
        dcache[2056] = 64'h822c0060809e8133;
        dcache[2057] = 64'h803f804a802b0029;
        dcache[2058] = 64'h01d000e501358053;
        dcache[2059] = 64'h0086802e809a8062;
        dcache[2060] = 64'h8239011a80e4815f;
        dcache[2061] = 64'h00d78035003e8022;
        dcache[2062] = 64'h00d900260170003d;
        dcache[2063] = 64'h00230072803d807c;
        dcache[2064] = 64'h81d700158112818b;
        dcache[2065] = 64'h016e0104804000dc;
        dcache[2066] = 64'h009e80d5016d0000;
        dcache[2067] = 64'h80f4003c812c80c8;
        dcache[2068] = 64'h80af006780488114;
        dcache[2069] = 64'h01fe00bc800400f7;
        dcache[2070] = 64'h8036803c015f005f;
        dcache[2071] = 64'h80d40098811b814d;
        dcache[2072] = 64'h0075803f80080015;
        dcache[2073] = 64'h010500a101340090;
        dcache[2074] = 64'h80770006010100c6;
        dcache[2075] = 64'h805300ca805480ee;
        dcache[2076] = 64'h0060801800580035;
        dcache[2077] = 64'h000b00fc0169800d;
        dcache[2078] = 64'h8008004b00870101;
        dcache[2079] = 64'h0076802c0032800e;
        dcache[2080] = 64'h8010806680040032;
        dcache[2081] = 64'h0045017c00e6000c;
        dcache[2082] = 64'h0077804e803a013e;
        dcache[2083] = 64'h00ec802700108027;
        dcache[2084] = 64'h8082807100120052;
        dcache[2085] = 64'h005101370088008e;
        dcache[2086] = 64'h800600d380130103;
        dcache[2087] = 64'h015e804780558022;
        dcache[2088] = 64'h80d480508020004b;
        dcache[2089] = 64'h00ae0114003e00d4;
        dcache[2090] = 64'h800600978008003f;
        dcache[2091] = 64'h00ce8016814c8098;
        dcache[2092] = 64'h80ec00820021002a;
        dcache[2093] = 64'h006b008a008e00bd;
        dcache[2094] = 64'h8034005300000076;
        dcache[2095] = 64'h0048000d80210024;
        dcache[2096] = 64'h80850068007b003c;
        dcache[2097] = 64'h0073004e005f8055;
        dcache[2098] = 64'h0013804a00630028;
        dcache[2099] = 64'h806b00a500398053;
        dcache[2100] = 64'h80a700ac00c50094;
        dcache[2101] = 64'h000f00ac010d806c;
        dcache[2102] = 64'h805080868083006a;
        dcache[2103] = 64'h003780a180228076;
        dcache[2104] = 64'h8203005501810064;
        dcache[2105] = 64'h80e900bb00b80016;
        dcache[2106] = 64'h8022804f80118063;
        dcache[2107] = 64'h00df80a680408016;
        dcache[2108] = 64'h829d005200db0022;
        dcache[2109] = 64'h8063012d00978100;
        dcache[2110] = 64'h010b810781368046;
        dcache[2111] = 64'h8043809f8076805e;
        dcache[2112] = 64'h8111800200d90074;
        dcache[2113] = 64'h007800a98012006a;
        dcache[2114] = 64'h00bc80a480f68160;
        dcache[2115] = 64'h808e80538006808d;
        dcache[2116] = 64'h8140806701bc0302;
        dcache[2117] = 64'h020101da016100b0;
        dcache[2118] = 64'h0059005780418207;
        dcache[2119] = 64'h004680af8238013c;
        dcache[2120] = 64'h8018803c00d680b1;
        dcache[2121] = 64'h0030808480de01ed;
        dcache[2122] = 64'h811e0008017080f1;
        dcache[2123] = 64'h010200e080bd804e;
        dcache[2124] = 64'h001980d801fb8072;
        dcache[2125] = 64'h007d01ce01dd0196;
        dcache[2126] = 64'h8176802000d78203;
        dcache[2127] = 64'h801a003e80bc0002;
        dcache[2128] = 64'h005f808700ac0046;
        dcache[2129] = 64'h8098005580a9001c;
        dcache[2130] = 64'h808200e70029001e;
        dcache[2131] = 64'h810300c1803580bd;
        dcache[2132] = 64'h010500de815c0067;
        dcache[2133] = 64'h8160801881678092;
        dcache[2134] = 64'h807e00ba0105814a;
        dcache[2135] = 64'h01ae800380f300a6;
        dcache[2136] = 64'h014c0196812500e6;
        dcache[2137] = 64'h006b814780728035;
        dcache[2138] = 64'h00950158006780ba;
        dcache[2139] = 64'h806500388065803f;
        dcache[2140] = 64'h8077019b00eb808b;
        dcache[2141] = 64'h00010086010e0094;
        dcache[2142] = 64'h80d3807482100135;
        dcache[2143] = 64'h00c18191800d8070;
        dcache[2144] = 64'h009001688037011f;
        dcache[2145] = 64'h801f00ae01c400fa;
        dcache[2146] = 64'h0060819d82060047;
        dcache[2147] = 64'h01018027009e0023;
        dcache[2148] = 64'h80d7014c002e8012;
        dcache[2149] = 64'h8045015400450084;
        dcache[2150] = 64'h008d814882e4007a;
        dcache[2151] = 64'h011f803e013f803c;
        dcache[2152] = 64'h8136015000470105;
        dcache[2153] = 64'h0091008780a500ce;
        dcache[2154] = 64'h0096807b82b60021;
        dcache[2155] = 64'h0008002400268042;
        dcache[2156] = 64'h820200d100c58027;
        dcache[2157] = 64'h001f00b2801d00ab;
        dcache[2158] = 64'h011f808380fc8090;
        dcache[2159] = 64'h002b80c980948030;
        dcache[2160] = 64'h82c2014b80438079;
        dcache[2161] = 64'h8027000e80b58017;
        dcache[2162] = 64'h010e805080e880d6;
        dcache[2163] = 64'h800a006e80a7800f;
        dcache[2164] = 64'h8273011a80288116;
        dcache[2165] = 64'h80080089813f0046;
        dcache[2166] = 64'h0155003e0046807d;
        dcache[2167] = 64'h8029800181728089;
        dcache[2168] = 64'h832c00d5802b80f7;
        dcache[2169] = 64'h005a00a780b58007;
        dcache[2170] = 64'h0118004b01798033;
        dcache[2171] = 64'h00238078814a8071;
        dcache[2172] = 64'h82e2009581e080f5;
        dcache[2173] = 64'h008b00d8809c006e;
        dcache[2174] = 64'h00b4805e01a6802f;
        dcache[2175] = 64'h80110012814c80df;
        dcache[2176] = 64'h8277004981bc8107;
        dcache[2177] = 64'h0079002280b00008;
        dcache[2178] = 64'h0064002201838011;
        dcache[2179] = 64'h0043802581810003;
        dcache[2180] = 64'h80c0006080f18039;
        dcache[2181] = 64'h00b200bd801c00ca;
        dcache[2182] = 64'h8012003f01788023;
        dcache[2183] = 64'h000c00068155803e;
        dcache[2184] = 64'h008c0062804c0067;
        dcache[2185] = 64'h008f011500880021;
        dcache[2186] = 64'h0026800d00d9008e;
        dcache[2187] = 64'h0046003b80bf8073;
        dcache[2188] = 64'h00460004005400c9;
        dcache[2189] = 64'h0036018000c90053;
        dcache[2190] = 64'h0049008e805700bd;
        dcache[2191] = 64'h80298031805f007b;
        dcache[2192] = 64'h80cc80d0012700ee;
        dcache[2193] = 64'h00a3013300b9001b;
        dcache[2194] = 64'h0025000e805d0097;
        dcache[2195] = 64'h8001808980a0800e;
        dcache[2196] = 64'h8124806500900046;
        dcache[2197] = 64'h001e019f8001007f;
        dcache[2198] = 64'h00a300208036008a;
        dcache[2199] = 64'h00b0803080350097;
        dcache[2200] = 64'h819c8099007e0071;
        dcache[2201] = 64'h800a015200288043;
        dcache[2202] = 64'h800b002e800500c1;
        dcache[2203] = 64'h8012802e800c0040;
        dcache[2204] = 64'h81750044005b007c;
        dcache[2205] = 64'h0022804800850027;
        dcache[2206] = 64'h801800560029008f;
        dcache[2207] = 64'h8043803a00550022;
        dcache[2208] = 64'h819d807e002a00d8;
        dcache[2209] = 64'h004700110021007b;
        dcache[2210] = 64'h003b8070001f8019;
        dcache[2211] = 64'h8001804a00a100ac;
        dcache[2212] = 64'h8185006900ef00f0;
        dcache[2213] = 64'h801e010a01220072;
        dcache[2214] = 64'h00cc812080e30057;
        dcache[2215] = 64'h0000810d00598071;
        dcache[2216] = 64'h834600630149006f;
        dcache[2217] = 64'h800f00f201030026;
        dcache[2218] = 64'h010f806380bb8097;
        dcache[2219] = 64'h802781b800388010;
        dcache[2220] = 64'h82ff007200dc0009;
        dcache[2221] = 64'h80a7007300190044;
        dcache[2222] = 64'h000a004880c88040;
        dcache[2223] = 64'h8119820d008f80c2;
        dcache[2224] = 64'h81af0006802200e9;
        dcache[2225] = 64'h8052805200ad0068;
        dcache[2226] = 64'h802800da80128162;
        dcache[2227] = 64'h8047800380240031;
        dcache[2228] = 64'h808a80d60140035b;
        dcache[2229] = 64'h0157015200850171;
        dcache[2230] = 64'h814800ad81708212;
        dcache[2231] = 64'h006c005c81b6005d;
        dcache[2232] = 64'h0119805a030d800d;
        dcache[2233] = 64'h0118021c01080230;
        dcache[2234] = 64'h001e80ed005482c5;
        dcache[2235] = 64'h00fd803e80140051;
        dcache[2236] = 64'h008780b8016e807d;
        dcache[2237] = 64'h0060017f018d011c;
        dcache[2238] = 64'h80cd8046011e820d;
        dcache[2239] = 64'h8080012f815d8069;
        dcache[2240] = 64'h001200360021004d;
        dcache[2241] = 64'h0020801f8013003b;
        dcache[2242] = 64'h8033002800088042;
        dcache[2243] = 64'h003a000780150006;
        dcache[2244] = 64'h002d0160802a80e4;
        dcache[2245] = 64'h80c4810e005c8029;
        dcache[2246] = 64'h00ff80678009803a;
        dcache[2247] = 64'h018d0133010b003c;
        dcache[2248] = 64'h010c0031809c0100;
        dcache[2249] = 64'h006000878032801e;
        dcache[2250] = 64'h00df80c682638065;
        dcache[2251] = 64'h805b803b002f0085;
        dcache[2252] = 64'h817100a100410022;
        dcache[2253] = 64'h806001cb00b801c2;
        dcache[2254] = 64'h805980bb83710069;
        dcache[2255] = 64'h00c881ba008000d5;
        dcache[2256] = 64'h81a200ad00e50159;
        dcache[2257] = 64'h80b500da00cb0151;
        dcache[2258] = 64'h003c80e383d48031;
        dcache[2259] = 64'h00d580d000cc012e;
        dcache[2260] = 64'h825f00e1800b0119;
        dcache[2261] = 64'h0042806a80670079;
        dcache[2262] = 64'h00cf80a48389803b;
        dcache[2263] = 64'h0113000b01150183;
        dcache[2264] = 64'h826200cf00970089;
        dcache[2265] = 64'h80a5003280be00a2;
        dcache[2266] = 64'h006880ad81648076;
        dcache[2267] = 64'h0051800d0094005e;
        dcache[2268] = 64'h838f00ae012000c8;
        dcache[2269] = 64'h80c9010f80890037;
        dcache[2270] = 64'h00f3000d808880f6;
        dcache[2271] = 64'h803b80e1800a0066;
        dcache[2272] = 64'h8290011a001d0073;
        dcache[2273] = 64'h80ac00818069002f;
        dcache[2274] = 64'h003a0067808480b7;
        dcache[2275] = 64'h001a002f80a90037;
        dcache[2276] = 64'h820a00e2802200bd;
        dcache[2277] = 64'h80b6015a80c40043;
        dcache[2278] = 64'h00a40032809b8008;
        dcache[2279] = 64'h8027806d80f08021;
        dcache[2280] = 64'h815900de8046804f;
        dcache[2281] = 64'h809500ca80b60001;
        dcache[2282] = 64'h014f0066005f8073;
        dcache[2283] = 64'h8045800b81158008;
        dcache[2284] = 64'h80eb005681460099;
        dcache[2285] = 64'h80aa00ef80aa0062;
        dcache[2286] = 64'h010900200076809e;
        dcache[2287] = 64'h00038057811f8017;
        dcache[2288] = 64'h806d8003814f006e;
        dcache[2289] = 64'h800600b580ed803e;
        dcache[2290] = 64'h00ad803901288095;
        dcache[2291] = 64'h801c007480f0007e;
        dcache[2292] = 64'h809700338075008b;
        dcache[2293] = 64'h8002006381260007;
        dcache[2294] = 64'h007a008f007c000a;
        dcache[2295] = 64'h0058802d803b00cc;
        dcache[2296] = 64'h0061004980340113;
        dcache[2297] = 64'h002100bc80b70032;
        dcache[2298] = 64'h000200c5009e015d;
        dcache[2299] = 64'h002f80b480d7007e;
        dcache[2300] = 64'h8023800d005200e3;
        dcache[2301] = 64'h005d00bf80fb8077;
        dcache[2302] = 64'h007e001b80500036;
        dcache[2303] = 64'h003d80aa805200ce;
        dcache[2304] = 64'h0005808200a50167;
        dcache[2305] = 64'h002f009f807c0049;
        dcache[2306] = 64'h8014006e808b007b;
        dcache[2307] = 64'h002a809b80160025;
        dcache[2308] = 64'h8005807700a300c7;
        dcache[2309] = 64'h005a00bb80658097;
        dcache[2310] = 64'h8044001580da00a8;
        dcache[2311] = 64'h801b8016008e007d;
        dcache[2312] = 64'h80e0803900bf00fe;
        dcache[2313] = 64'h0012011c00658006;
        dcache[2314] = 64'h001f007d8022004d;
        dcache[2315] = 64'h80b98083802d007c;
        dcache[2316] = 64'h81cc804e00970175;
        dcache[2317] = 64'h800380110021001a;
        dcache[2318] = 64'h802e80230021802c;
        dcache[2319] = 64'h803880c7004e0038;
        dcache[2320] = 64'h81a680bf010400eb;
        dcache[2321] = 64'h804800c081170055;
        dcache[2322] = 64'h80168079806d005d;
        dcache[2323] = 64'h803f811300900097;
        dcache[2324] = 64'h815a0027008f012c;
        dcache[2325] = 64'h005d00db80460002;
        dcache[2326] = 64'h00be811d80e68047;
        dcache[2327] = 64'h808a817600f30099;
        dcache[2328] = 64'h82540092007100f8;
        dcache[2329] = 64'h80428028001d8072;
        dcache[2330] = 64'h006380c08111804c;
        dcache[2331] = 64'h80ae810401300116;
        dcache[2332] = 64'h82980125006700da;
        dcache[2333] = 64'h00240007000e0093;
        dcache[2334] = 64'h8003804281098085;
        dcache[2335] = 64'h80d881c1007f009d;
        dcache[2336] = 64'h81a88069801f0040;
        dcache[2337] = 64'h0117810900dc000d;
        dcache[2338] = 64'h80e6005d007a8181;
        dcache[2339] = 64'h00318024007a800f;
        dcache[2340] = 64'h810380dc80590242;
        dcache[2341] = 64'h01c4808e006e0117;
        dcache[2342] = 64'h820d017f808c811a;
        dcache[2343] = 64'h801b800c002c8029;
        dcache[2344] = 64'h000580ce01590080;
        dcache[2345] = 64'h000101df80260128;
        dcache[2346] = 64'h800e00640109827e;
        dcache[2347] = 64'h805b003a812280a0;
        dcache[2348] = 64'h801f804c00d6000a;
        dcache[2349] = 64'h813a0141807d0007;
        dcache[2350] = 64'h815700fd006f0091;
        dcache[2351] = 64'h8087015d801880e6;
        dcache[2352] = 64'h001a80d200a60046;
        dcache[2353] = 64'h80df00cd003c007d;
        dcache[2354] = 64'h8109010a007d808e;
        dcache[2355] = 64'h8141010c80bc8093;
        dcache[2356] = 64'h80270023019b80d8;
        dcache[2357] = 64'h801500f6007b00e7;
        dcache[2358] = 64'h802e007d80f8006f;
        dcache[2359] = 64'h013381528026802d;
        dcache[2360] = 64'h813880390217001c;
        dcache[2361] = 64'h80b6023c8093015f;
        dcache[2362] = 64'h0014807381d70011;
        dcache[2363] = 64'h803482b00091026c;
        dcache[2364] = 64'h820481430066012e;
        dcache[2365] = 64'h806e027180230168;
        dcache[2366] = 64'h0043807d82878001;
        dcache[2367] = 64'h807280fd0069016b;
        dcache[2368] = 64'h822280450120013a;
        dcache[2369] = 64'h8049004c00090013;
        dcache[2370] = 64'h8008800582338005;
        dcache[2371] = 64'h808c806300e80001;
        dcache[2372] = 64'h82ac803c00750100;
        dcache[2373] = 64'h0027806f002a006a;
        dcache[2374] = 64'h806d801f818980ad;
        dcache[2375] = 64'h809e007b800d805c;
        dcache[2376] = 64'h82c9002200be00e2;
        dcache[2377] = 64'h805880a180c28082;
        dcache[2378] = 64'h8030801680a780cc;
        dcache[2379] = 64'h8021003100bb004e;
        dcache[2380] = 64'h82360021007e00cc;
        dcache[2381] = 64'h80c5001b80738090;
        dcache[2382] = 64'h008300d680838059;
        dcache[2383] = 64'h8054800200c30044;
        dcache[2384] = 64'h80818007006a0143;
        dcache[2385] = 64'h8044001e809a80a0;
        dcache[2386] = 64'h0016007580a10052;
        dcache[2387] = 64'h0006802380240051;
        dcache[2388] = 64'h8023806180040112;
        dcache[2389] = 64'h001d004c80e88053;
        dcache[2390] = 64'h0162800d8041805a;
        dcache[2391] = 64'h805e80588084000e;
        dcache[2392] = 64'h8000001c800f0105;
        dcache[2393] = 64'h8021001480df0056;
        dcache[2394] = 64'h010400b280058017;
        dcache[2395] = 64'h8007804780820082;
        dcache[2396] = 64'h802600a380880105;
        dcache[2397] = 64'h000300158101801a;
        dcache[2398] = 64'h00f4002580158013;
        dcache[2399] = 64'h806b804b803b0102;
        dcache[2400] = 64'h808e007c80e80136;
        dcache[2401] = 64'h8066006d80998039;
        dcache[2402] = 64'h00d3008c003b001f;
        dcache[2403] = 64'h8025808f803300fc;
        dcache[2404] = 64'h80510060806d00f3;
        dcache[2405] = 64'h00a900a28152000e;
        dcache[2406] = 64'h00fb00c60080009a;
        dcache[2407] = 64'h803880de804a00f6;
        dcache[2408] = 64'h806600a780460184;
        dcache[2409] = 64'h801600408198805a;
        dcache[2410] = 64'h0069007e00d700cc;
        dcache[2411] = 64'h808880a7804b0115;
        dcache[2412] = 64'h0009002f000d0134;
        dcache[2413] = 64'h8018004482008088;
        dcache[2414] = 64'h0059004800430067;
        dcache[2415] = 64'h80328067805600df;
        dcache[2416] = 64'h80368001004400ea;
        dcache[2417] = 64'h0052004581080035;
        dcache[2418] = 64'h0011007a80360053;
        dcache[2419] = 64'h0081812e808e006e;
        dcache[2420] = 64'h805b000d010300a1;
        dcache[2421] = 64'h011b00a581c90016;
        dcache[2422] = 64'h006a003a80a00005;
        dcache[2423] = 64'h8080806f806a0090;
        dcache[2424] = 64'h805e8048008f00e9;
        dcache[2425] = 64'h0021006f80f6001d;
        dcache[2426] = 64'h8041802180050008;
        dcache[2427] = 64'h80a380ff80cc0021;
        dcache[2428] = 64'h80e78036005900f2;
        dcache[2429] = 64'h00a100148125008f;
        dcache[2430] = 64'h803f807280668062;
        dcache[2431] = 64'h80fc810a804e00be;
        dcache[2432] = 64'h812580cc00120115;
        dcache[2433] = 64'h009280638193002a;
        dcache[2434] = 64'h806f8007804b8021;
        dcache[2435] = 64'h8158809600470068;
        dcache[2436] = 64'h810780c400390168;
        dcache[2437] = 64'h001c8004002700dd;
        dcache[2438] = 64'h805080bb807d8072;
        dcache[2439] = 64'h816e80dc004a0111;
        dcache[2440] = 64'h80b400fb0036017e;
        dcache[2441] = 64'h007a000880230099;
        dcache[2442] = 64'h012781b281950013;
        dcache[2443] = 64'h810c814e00a201b1;
        dcache[2444] = 64'h8105004180340191;
        dcache[2445] = 64'h017300e1803c0099;
        dcache[2446] = 64'h006881cc80be812c;
        dcache[2447] = 64'h804e815a010d0200;
        dcache[2448] = 64'h805c80df00260235;
        dcache[2449] = 64'h01c4805d804c8011;
        dcache[2450] = 64'h82150082805581e4;
        dcache[2451] = 64'h8112000a002a804e;
        dcache[2452] = 64'h8090818d005e024a;
        dcache[2453] = 64'h00ab002381250071;
        dcache[2454] = 64'h81da00b200ad8146;
        dcache[2455] = 64'h807f004c00038044;
        dcache[2456] = 64'h81178029812500f4;
        dcache[2457] = 64'h8012018a003b00b9;
        dcache[2458] = 64'h019681640023817b;
        dcache[2459] = 64'h019a8000802d00bf;
        dcache[2460] = 64'h00480028000e8039;
        dcache[2461] = 64'h8067801980160029;
        dcache[2462] = 64'h004b800e802a004e;
        dcache[2463] = 64'h0072001e8055005d;
        dcache[2464] = 64'h002380a7008a0008;
        dcache[2465] = 64'h8124009f00340012;
        dcache[2466] = 64'h80ad00b500c0805f;
        dcache[2467] = 64'h8133012e80e88100;
        dcache[2468] = 64'h805f0007007c80ec;
        dcache[2469] = 64'h80c80078002c0044;
        dcache[2470] = 64'h81250129003a011a;
        dcache[2471] = 64'h80410078801e8121;
        dcache[2472] = 64'h81900008022f8007;
        dcache[2473] = 64'h005001d68033018a;
        dcache[2474] = 64'h006b801481bc801e;
        dcache[2475] = 64'h005c82a70017020c;
        dcache[2476] = 64'h823e803201d40172;
        dcache[2477] = 64'h001b020f0008009c;
        dcache[2478] = 64'h0024000d82b60097;
        dcache[2479] = 64'h807481100095016b;
        dcache[2480] = 64'h820e000400ed016f;
        dcache[2481] = 64'h00a7014180200147;
        dcache[2482] = 64'h803f0008815e807a;
        dcache[2483] = 64'h8154802201060015;
        dcache[2484] = 64'h82bd809d02370079;
        dcache[2485] = 64'h0039003680aa0195;
        dcache[2486] = 64'h807c0048006181cd;
        dcache[2487] = 64'h80c9800b81398016;
        dcache[2488] = 64'h81c88029016d0040;
        dcache[2489] = 64'h806080b0809a804b;
        dcache[2490] = 64'h8034806180ac8173;
        dcache[2491] = 64'h80200107803700bc;
        dcache[2492] = 64'h800b003d01260106;
        dcache[2493] = 64'h8047001f804d8039;
        dcache[2494] = 64'h0015807d8081809a;
        dcache[2495] = 64'h00510036800400c0;
        dcache[2496] = 64'h0146807f0030017a;
        dcache[2497] = 64'h0025804a80780011;
        dcache[2498] = 64'h0055800a811580dc;
        dcache[2499] = 64'h0099802d803d0148;
        dcache[2500] = 64'h00cb0019002200f1;
        dcache[2501] = 64'h00530029805a8069;
        dcache[2502] = 64'h0054000e8068802f;
        dcache[2503] = 64'h003d802c80e90169;
        dcache[2504] = 64'h007580140016004e;
        dcache[2505] = 64'h0021803580318031;
        dcache[2506] = 64'h00d7001f8074005f;
        dcache[2507] = 64'h00328041808e0067;
        dcache[2508] = 64'h806b0083806d0046;
        dcache[2509] = 64'h8006803a8192806e;
        dcache[2510] = 64'h00f68012809500a4;
        dcache[2511] = 64'h000d000d802600ef;
        dcache[2512] = 64'h0017007e80e100e6;
        dcache[2513] = 64'h006a805f80e380bc;
        dcache[2514] = 64'h013d0020004400bb;
        dcache[2515] = 64'h001d807280270110;
        dcache[2516] = 64'h0011801280da0096;
        dcache[2517] = 64'h801c0007812a003f;
        dcache[2518] = 64'h0162004e00190085;
        dcache[2519] = 64'h804f8011003c0120;
        dcache[2520] = 64'h003c003b000c00c4;
        dcache[2521] = 64'h804780a481bd000f;
        dcache[2522] = 64'h00c500ae007a00f3;
        dcache[2523] = 64'h00180018001100b0;
        dcache[2524] = 64'h007100038090010d;
        dcache[2525] = 64'h807e801b819e804c;
        dcache[2526] = 64'h0069003a00c00163;
        dcache[2527] = 64'h804680af80760108;
        dcache[2528] = 64'h00278004001600bd;
        dcache[2529] = 64'h8046804f81918001;
        dcache[2530] = 64'h00268001001200d5;
        dcache[2531] = 64'h0013807f0036010f;
        dcache[2532] = 64'h001b8046007d0039;
        dcache[2533] = 64'h0015000681fd009b;
        dcache[2534] = 64'h80b3800e80a00057;
        dcache[2535] = 64'h805e8075806b00fd;
        dcache[2536] = 64'h80308016007b00d2;
        dcache[2537] = 64'h801b80b68117004c;
        dcache[2538] = 64'h805c80b180ac0009;
        dcache[2539] = 64'h812880b3806c00e6;
        dcache[2540] = 64'h0012001e004600b2;
        dcache[2541] = 64'h004700aa81fa006d;
        dcache[2542] = 64'h8056817881300062;
        dcache[2543] = 64'h811d80bf805000cd;
        dcache[2544] = 64'h8104817f00ab00fa;
        dcache[2545] = 64'h0048803380ff0042;
        dcache[2546] = 64'h8098801c80b2003c;
        dcache[2547] = 64'h812b81378020006e;
        dcache[2548] = 64'h802f818b00a8015b;
        dcache[2549] = 64'h00a6003680450094;
        dcache[2550] = 64'h000c818680840052;
        dcache[2551] = 64'h814481fb802b0090;
        dcache[2552] = 64'h0055008f008800ea;
        dcache[2553] = 64'h004480b380320006;
        dcache[2554] = 64'h0063817080b10034;
        dcache[2555] = 64'h007c80ef01460192;
        dcache[2556] = 64'h808e8025000f01bd;
        dcache[2557] = 64'h00b380b18059803b;
        dcache[2558] = 64'h80718055802480c6;
        dcache[2559] = 64'h000300b2013c0214;
        dcache[2560] = 64'h80078138002f00e2;
        dcache[2561] = 64'h025d808f8016803e;
        dcache[2562] = 64'h80d80085006081bd;
        dcache[2563] = 64'h808f00940098008d;
        dcache[2564] = 64'h805481db00a7021f;
        dcache[2565] = 64'h8013001b80ea801e;
        dcache[2566] = 64'h81390110006f8113;
        dcache[2567] = 64'h80fd005c80258064;
        dcache[2568] = 64'h0047806980a30120;
        dcache[2569] = 64'h81f80074810e80a8;
        dcache[2570] = 64'h80e800bb80b300b4;
        dcache[2571] = 64'h81cb01cd008480c7;
        dcache[2572] = 64'h803580618070004f;
        dcache[2573] = 64'h802480570027000e;
        dcache[2574] = 64'h00148039001d0052;
        dcache[2575] = 64'h006f804380510002;
        dcache[2576] = 64'h801b003e003c002b;
        dcache[2577] = 64'h803a002d803e0041;
        dcache[2578] = 64'h0010000880258014;
        dcache[2579] = 64'h80190052000a0007;
        dcache[2580] = 64'h803f0050802e0015;
        dcache[2581] = 64'h001e0022003a0056;
        dcache[2582] = 64'h0025802d80158020;
        dcache[2583] = 64'h003600338036802e;
        dcache[2584] = 64'h81da01c001ea0003;
        dcache[2585] = 64'h80f502010064006c;
        dcache[2586] = 64'h805000fe81a8011c;
        dcache[2587] = 64'h8042829000b7024e;
        dcache[2588] = 64'h81600138011e00e2;
        dcache[2589] = 64'h806001890023003e;
        dcache[2590] = 64'h807d009d835e0255;
        dcache[2591] = 64'h0101823002630196;
        dcache[2592] = 64'h818801e0802b014e;
        dcache[2593] = 64'h0071008a81330000;
        dcache[2594] = 64'h8027807c810e0040;
        dcache[2595] = 64'h005380d1016900b7;
        dcache[2596] = 64'h80fb0070005e010c;
        dcache[2597] = 64'h0064001580f9008c;
        dcache[2598] = 64'h80f7003680ef8098;
        dcache[2599] = 64'h005e001780840083;
        dcache[2600] = 64'h8030004880590057;
        dcache[2601] = 64'h806980c8808500af;
        dcache[2602] = 64'h80ea812581158050;
        dcache[2603] = 64'h00df803880a0006f;
        dcache[2604] = 64'h0046001100cb0025;
        dcache[2605] = 64'h80ca80ac80470097;
        dcache[2606] = 64'h8051812000018032;
        dcache[2607] = 64'h017e001880420153;
        dcache[2608] = 64'h8011803a00eb009b;
        dcache[2609] = 64'h8019804a808a8025;
        dcache[2610] = 64'h006380f381080029;
        dcache[2611] = 64'h004c008f0115014a;
        dcache[2612] = 64'h0092806100db0047;
        dcache[2613] = 64'h8029004e80c78054;
        dcache[2614] = 64'h004480cb80548023;
        dcache[2615] = 64'h000f0056805a0170;
        dcache[2616] = 64'h803f0067002b00a9;
        dcache[2617] = 64'h8056002e80468087;
        dcache[2618] = 64'h000180f7807b0027;
        dcache[2619] = 64'h00e200f1009f0189;
        dcache[2620] = 64'h8081008700370092;
        dcache[2621] = 64'h80510047803f0052;
        dcache[2622] = 64'h004480508042007f;
        dcache[2623] = 64'h009a0035007f01bf;
        dcache[2624] = 64'h0024806b002f0083;
        dcache[2625] = 64'h801400418074006b;
        dcache[2626] = 64'h0092000000a3803b;
        dcache[2627] = 64'h000600f5800e014e;
        dcache[2628] = 64'h8030003a0080006e;
        dcache[2629] = 64'h80c2800c813100a0;
        dcache[2630] = 64'h008a802100630079;
        dcache[2631] = 64'h802500670081012a;
        dcache[2632] = 64'h00a38047809000c4;
        dcache[2633] = 64'h8076805c80c9803c;
        dcache[2634] = 64'h007980b1004900a2;
        dcache[2635] = 64'h800d0069004a00f7;
        dcache[2636] = 64'h0078001c800500b0;
        dcache[2637] = 64'h807f8027815c8032;
        dcache[2638] = 64'h0088803200d600cf;
        dcache[2639] = 64'h807b0010002200f0;
        dcache[2640] = 64'h00bf000a0015007a;
        dcache[2641] = 64'h0040806a815c802f;
        dcache[2642] = 64'h002680830035006a;
        dcache[2643] = 64'h80b6004900a60100;
        dcache[2644] = 64'h0045804800e800bc;
        dcache[2645] = 64'h809580e881b68054;
        dcache[2646] = 64'h806880c0005600de;
        dcache[2647] = 64'h810880220006017a;
        dcache[2648] = 64'h000c807b016c0018;
        dcache[2649] = 64'h006680c581368002;
        dcache[2650] = 64'h00328115801e0097;
        dcache[2651] = 64'h8154818980070094;
        dcache[2652] = 64'h0046806b00b7002c;
        dcache[2653] = 64'h009e807880f9000b;
        dcache[2654] = 64'h002a80fc802a800d;
        dcache[2655] = 64'h8101813780e2010e;
        dcache[2656] = 64'h001180e4015000d9;
        dcache[2657] = 64'h0168801b80ee8081;
        dcache[2658] = 64'h805f804280580081;
        dcache[2659] = 64'h80e8816c801200be;
        dcache[2660] = 64'h00b7812c01050087;
        dcache[2661] = 64'h022a808280bb8072;
        dcache[2662] = 64'h001a81378000003c;
        dcache[2663] = 64'h80e181a500b300f7;
        dcache[2664] = 64'h80c180f401600112;
        dcache[2665] = 64'h01b581330029005d;
        dcache[2666] = 64'h00990081000a812d;
        dcache[2667] = 64'h0034813f014f0297;
        dcache[2668] = 64'h81b280b1013400f3;
        dcache[2669] = 64'h029980b88054803b;
        dcache[2670] = 64'h004f005f005180db;
        dcache[2671] = 64'h80538072032e0266;
        dcache[2672] = 64'h817e807100560109;
        dcache[2673] = 64'h020e80e9005f00db;
        dcache[2674] = 64'h81180122006f80ee;
        dcache[2675] = 64'h00ee0030009c01b8;
        dcache[2676] = 64'h801f8081003c0172;
        dcache[2677] = 64'h0124804d809a8049;
        dcache[2678] = 64'h805c0004001080ad;
        dcache[2679] = 64'h809f0087800c00bc;
        dcache[2680] = 64'h012c808e806201e8;
        dcache[2681] = 64'h8131018e0048005e;
        dcache[2682] = 64'h81ab0128804b0102;
        dcache[2683] = 64'h82a7013f808f8196;
        dcache[2684] = 64'h0042803f803f001f;
        dcache[2685] = 64'h803a001d80200022;
        dcache[2686] = 64'h0044804b801c001a;
        dcache[2687] = 64'h0044003e001a0050;
        dcache[2688] = 64'h80098028001a0038;
        dcache[2689] = 64'h80530015802b0041;
        dcache[2690] = 64'h0004002d0006001d;
        dcache[2691] = 64'h8039801480048017;
        dcache[2692] = 64'h002d000b00050022;
        dcache[2693] = 64'h8047000800400005;
        dcache[2694] = 64'h000b00140049001f;
        dcache[2695] = 64'h0049004e80070012;
        dcache[2696] = 64'h00dc8027010680e1;
        dcache[2697] = 64'h003f011080e5010f;
        dcache[2698] = 64'h0017805800468055;
        dcache[2699] = 64'h00c4815380a7805d;
        dcache[2700] = 64'h000d028580dc80fa;
        dcache[2701] = 64'h81e7804f81680071;
        dcache[2702] = 64'h81de019381a40276;
        dcache[2703] = 64'h01f3811401a30055;
        dcache[2704] = 64'h80fc00748146801e;
        dcache[2705] = 64'h81b581f4008000bc;
        dcache[2706] = 64'h811700be00310217;
        dcache[2707] = 64'h03f1819500a8001a;
        dcache[2708] = 64'h8011002f812d00bf;
        dcache[2709] = 64'h808581bd006d8053;
        dcache[2710] = 64'h8111800b00920135;
        dcache[2711] = 64'h027d005d80a78145;
        dcache[2712] = 64'h809200e7816f0126;
        dcache[2713] = 64'h80d0816080698020;
        dcache[2714] = 64'h811180fb005a01a0;
        dcache[2715] = 64'h01248047002b8051;
        dcache[2716] = 64'h80a9004380ad0114;
        dcache[2717] = 64'h806781d90043001d;
        dcache[2718] = 64'h81008119002c013f;
        dcache[2719] = 64'h00948032001e80a8;
        dcache[2720] = 64'h80710084809100c1;
        dcache[2721] = 64'h80478112808d0079;
        dcache[2722] = 64'h003980be001100d8;
        dcache[2723] = 64'h00340041009800bc;
        dcache[2724] = 64'h80650048806d0138;
        dcache[2725] = 64'h800d803e8082008c;
        dcache[2726] = 64'h000c80b180af00fd;
        dcache[2727] = 64'h803500d4003c010a;
        dcache[2728] = 64'h80fc004880650007;
        dcache[2729] = 64'h805180b98036001e;
        dcache[2730] = 64'h001e800580030196;
        dcache[2731] = 64'h0067004d0082009d;
        dcache[2732] = 64'h8046004b008e8001;
        dcache[2733] = 64'h005f801080cb803d;
        dcache[2734] = 64'h001980be00010132;
        dcache[2735] = 64'h005200cc010900a9;
        dcache[2736] = 64'h80f0005580230068;
        dcache[2737] = 64'h802d80a280c10063;
        dcache[2738] = 64'h00d2809f00150072;
        dcache[2739] = 64'h803800b400f901ad;
        dcache[2740] = 64'h801a009f809e8017;
        dcache[2741] = 64'h80a7805c80aa802d;
        dcache[2742] = 64'h009c805480b9009c;
        dcache[2743] = 64'h806300f801140122;
        dcache[2744] = 64'h800600dd80120099;
        dcache[2745] = 64'h808b000380e6005a;
        dcache[2746] = 64'h00ab80ff807f0038;
        dcache[2747] = 64'h80818006005e01b6;
        dcache[2748] = 64'h000300b600140069;
        dcache[2749] = 64'h807c807180eb809d;
        dcache[2750] = 64'h009b005000410088;
        dcache[2751] = 64'h8074001c007601e7;
        dcache[2752] = 64'h0072005680250004;
        dcache[2753] = 64'h000880a380fe80a6;
        dcache[2754] = 64'h00b68070003b0125;
        dcache[2755] = 64'h80c080e501b8017b;
        dcache[2756] = 64'h005d8025804900f8;
        dcache[2757] = 64'h80398074806c000e;
        dcache[2758] = 64'h80d0003680570055;
        dcache[2759] = 64'h804880ef8006016f;
        dcache[2760] = 64'h801e801800a40132;
        dcache[2761] = 64'h00e980d6800d8145;
        dcache[2762] = 64'h8025003a805b8043;
        dcache[2763] = 64'h815c80d2004c020f;
        dcache[2764] = 64'h801f807b00c9001c;
        dcache[2765] = 64'h011f805b801a8125;
        dcache[2766] = 64'h8134801f013b8061;
        dcache[2767] = 64'h8101805600d60175;
        dcache[2768] = 64'h001c8084000a007d;
        dcache[2769] = 64'h01768093002080cd;
        dcache[2770] = 64'h81fe00a200490077;
        dcache[2771] = 64'h002b809200f9015a;
        dcache[2772] = 64'h009b807900890073;
        dcache[2773] = 64'h01e000270024807c;
        dcache[2774] = 64'h826f00170040804f;
        dcache[2775] = 64'h006d818300350210;
        dcache[2776] = 64'h80898056800200bd;
        dcache[2777] = 64'h023480b801008005;
        dcache[2778] = 64'h8167804380f28010;
        dcache[2779] = 64'h0044806b00d60117;
        dcache[2780] = 64'h817d803200c3001c;
        dcache[2781] = 64'h023f804b00630033;
        dcache[2782] = 64'h8053006c8026003c;
        dcache[2783] = 64'h8063005803480098;
        dcache[2784] = 64'h80be800f0016010a;
        dcache[2785] = 64'h01cc00b600430269;
        dcache[2786] = 64'h810d00ae0015820f;
        dcache[2787] = 64'h012c8057001d026f;
        dcache[2788] = 64'h00d380f301d300f6;
        dcache[2789] = 64'h01f7018b013700bc;
        dcache[2790] = 64'h00d5819c00028189;
        dcache[2791] = 64'h003e80c1826b00e3;
        dcache[2792] = 64'h803280e300e80143;
        dcache[2793] = 64'h80a300d7003f0089;
        dcache[2794] = 64'h804f000a000680b7;
        dcache[2795] = 64'h804e808d81778006;
        dcache[2796] = 64'h8016800b000a0043;
        dcache[2797] = 64'h0051803d002a8020;
        dcache[2798] = 64'h8046004d00560013;
        dcache[2799] = 64'h000e803700438011;
        dcache[2800] = 64'h001d005700210037;
        dcache[2801] = 64'h0017001f00340031;
        dcache[2802] = 64'h003880400005801c;
        dcache[2803] = 64'h001f80548035802b;
        dcache[2804] = 64'h0046801800168007;
        dcache[2805] = 64'h8014802980298041;
        dcache[2806] = 64'h0056802380060052;
        dcache[2807] = 64'h8023002f8045800f;
        dcache[2808] = 64'h8120805f00a70056;
        dcache[2809] = 64'h8012003a00f1003b;
        dcache[2810] = 64'h812e018d81160159;
        dcache[2811] = 64'h00420006010c8059;
        dcache[2812] = 64'h0091808b815a00e1;
        dcache[2813] = 64'h014080ec80f20093;
        dcache[2814] = 64'h812c80b7004a80d3;
        dcache[2815] = 64'h8039014d806681d0;
        dcache[2816] = 64'h80ef8070825d80cb;
        dcache[2817] = 64'h00c581d70107005d;
        dcache[2818] = 64'h811a808e0155002d;
        dcache[2819] = 64'h0177008180c7806f;
        dcache[2820] = 64'h8133003582af80ca;
        dcache[2821] = 64'h802581ea022d8009;
        dcache[2822] = 64'h81ba015c002901a3;
        dcache[2823] = 64'h02998115001580b7;
        dcache[2824] = 64'h804601fa823d8003;
        dcache[2825] = 64'h801281b900298030;
        dcache[2826] = 64'h812d003e0096015e;
        dcache[2827] = 64'h00da818e0078801f;
        dcache[2828] = 64'h80ea01578207805c;
        dcache[2829] = 64'h807b8301004a00c4;
        dcache[2830] = 64'h819300a9010f012a;
        dcache[2831] = 64'h015881000075809a;
        dcache[2832] = 64'h8059012c80898091;
        dcache[2833] = 64'h80f682b3008b0174;
        dcache[2834] = 64'h8181019801050203;
        dcache[2835] = 64'h020480e200108014;
        dcache[2836] = 64'h001a01da810b006b;
        dcache[2837] = 64'h80738107003c0146;
        dcache[2838] = 64'h817f0123007601b5;
        dcache[2839] = 64'h0134003a008900ae;
        dcache[2840] = 64'h8088021481588056;
        dcache[2841] = 64'h01768108006e00f1;
        dcache[2842] = 64'h8043801a00210276;
        dcache[2843] = 64'h01b6808f02090057;
        dcache[2844] = 64'h00170209818e0025;
        dcache[2845] = 64'h011a815a004b005c;
        dcache[2846] = 64'h80c3002b007500f8;
        dcache[2847] = 64'h01260006018b0139;
        dcache[2848] = 64'h804d02c780990009;
        dcache[2849] = 64'h8004811e0024012c;
        dcache[2850] = 64'h81390158800400b8;
        dcache[2851] = 64'h00b9808600d00108;
        dcache[2852] = 64'h802c022080728053;
        dcache[2853] = 64'h0032818000578047;
        dcache[2854] = 64'h812900c88065010e;
        dcache[2855] = 64'h0029802901c400ab;
        dcache[2856] = 64'h8038018a003180be;
        dcache[2857] = 64'h019c819700230000;
        dcache[2858] = 64'h80d6008b00a70036;
        dcache[2859] = 64'h0033805c01470038;
        dcache[2860] = 64'h00ae01ca80578001;
        dcache[2861] = 64'h014d814b803100e0;
        dcache[2862] = 64'h814800428099807f;
        dcache[2863] = 64'h8051002001af01ee;
        dcache[2864] = 64'h8009024880558069;
        dcache[2865] = 64'h8001814a000b0030;
        dcache[2866] = 64'h815b012780648014;
        dcache[2867] = 64'h008d8069025a0168;
        dcache[2868] = 64'h003d025200258067;
        dcache[2869] = 64'h00d9817600478110;
        dcache[2870] = 64'h81d600e7001e0030;
        dcache[2871] = 64'h0025802e01c30093;
        dcache[2872] = 64'h000601a780c90023;
        dcache[2873] = 64'h009180d38027817e;
        dcache[2874] = 64'h81f4012f806800a5;
        dcache[2875] = 64'h8094802801b500b1;
        dcache[2876] = 64'h81350278812400cf;
        dcache[2877] = 64'h8107812b80748165;
        dcache[2878] = 64'h823a0176807f0147;
        dcache[2879] = 64'h007f803f01e6023a;
        dcache[2880] = 64'h8074001980338061;
        dcache[2881] = 64'h00c480e0002a812a;
        dcache[2882] = 64'h81f0017d801f0052;
        dcache[2883] = 64'h0017002e018b0161;
        dcache[2884] = 64'h0055000780538039;
        dcache[2885] = 64'h008a813580848184;
        dcache[2886] = 64'h82b401fa80ad0083;
        dcache[2887] = 64'h006f013c00e100fd;
        dcache[2888] = 64'h003e00e4822d01e0;
        dcache[2889] = 64'h804a8042811281d1;
        dcache[2890] = 64'h825b011b80ac0064;
        dcache[2891] = 64'h0012014000d50088;
        dcache[2892] = 64'h8076002d816e0156;
        dcache[2893] = 64'h8069007d804c805f;
        dcache[2894] = 64'h821800b880910222;
        dcache[2895] = 64'h8174014902e00008;
        dcache[2896] = 64'h80830111819f0144;
        dcache[2897] = 64'h8279004f80bf0087;
        dcache[2898] = 64'h82a2024c80320095;
        dcache[2899] = 64'h80ad00c702cd010d;
        dcache[2900] = 64'h0059807780260036;
        dcache[2901] = 64'h00fc809801080099;
        dcache[2902] = 64'h8088005580900063;
        dcache[2903] = 64'h01088100803d8075;
        dcache[2904] = 64'h801d800000010080;
        dcache[2905] = 64'h00730082004b008e;
        dcache[2906] = 64'h00b580a680638085;
        dcache[2907] = 64'h803880de806a00ce;
        dcache[2908] = 64'h0004801d001c000b;
        dcache[2909] = 64'h80520046804d8050;
        dcache[2910] = 64'h0052002c00150015;
        dcache[2911] = 64'h801b80420050804e;
        dcache[2912] = 64'h8051001300540031;
        dcache[2913] = 64'h802e000600420010;
        dcache[2914] = 64'h0045004400030044;
        dcache[2915] = 64'h8035800e00260028;
        dcache[2916] = 64'h0031000f801a8051;
        dcache[2917] = 64'h80100014803e0003;
        dcache[2918] = 64'h801b000e80348039;
        dcache[2919] = 64'h801d0006002b0049;
        dcache[2920] = 64'h8011804e80468047;
        dcache[2921] = 64'h80208053800a8003;
        dcache[2922] = 64'h805680130047001b;
        dcache[2923] = 64'h801d002a003d8037;
        dcache[2924] = 64'h001b80d400b5002a;
        dcache[2925] = 64'h007a80d100ec0034;
        dcache[2926] = 64'h005e00dc004100a5;
        dcache[2927] = 64'h00738008006d8040;
        dcache[2928] = 64'h8150817c00430035;
        dcache[2929] = 64'h019581570233807c;
        dcache[2930] = 64'h00ee001e80e50172;
        dcache[2931] = 64'h8067801201d9007e;
        dcache[2932] = 64'h819f8161818e807a;
        dcache[2933] = 64'h00e6815c02ee8159;
        dcache[2934] = 64'h0000007f80fd020a;
        dcache[2935] = 64'h001c80ef01aa807b;
        dcache[2936] = 64'h81348107827080c2;
        dcache[2937] = 64'h00d281ba02a68127;
        dcache[2938] = 64'h8055009e800101d1;
        dcache[2939] = 64'h011381ca017480f1;
        dcache[2940] = 64'h81640026801e8132;
        dcache[2941] = 64'h006482c701e80039;
        dcache[2942] = 64'h80fe02a301b4005d;
        dcache[2943] = 64'h026d821001128092;
        dcache[2944] = 64'h0040006200fd8248;
        dcache[2945] = 64'h00ac823400f9009f;
        dcache[2946] = 64'h80a0017d01c7006d;
        dcache[2947] = 64'h0298818300330055;
        dcache[2948] = 64'h00138029008081d4;
        dcache[2949] = 64'h008382c401670060;
        dcache[2950] = 64'h819d029d019e002d;
        dcache[2951] = 64'h0310811d0028000a;
        dcache[2952] = 64'h8017802400b28095;
        dcache[2953] = 64'h002981f801110059;
        dcache[2954] = 64'h82120226007700c7;
        dcache[2955] = 64'h02ca827100c000b8;
        dcache[2956] = 64'h808a006700478147;
        dcache[2957] = 64'h005a828c006e8053;
        dcache[2958] = 64'h8148023d002b00ae;
        dcache[2959] = 64'h01fb80fd012f016f;
        dcache[2960] = 64'h80810026002f822d;
        dcache[2961] = 64'h012a82f4007a80d5;
        dcache[2962] = 64'h00130281801d006b;
        dcache[2963] = 64'h01f0809301f50114;
        dcache[2964] = 64'h801400cf80fa8148;
        dcache[2965] = 64'h004282c1802c80f3;
        dcache[2966] = 64'h811003770005008c;
        dcache[2967] = 64'h02738044015e01a0;
        dcache[2968] = 64'h80648038000880c8;
        dcache[2969] = 64'h00c1843a01548033;
        dcache[2970] = 64'h818e045d000800b3;
        dcache[2971] = 64'h035980fa0173800b;
        dcache[2972] = 64'h00600038805580e1;
        dcache[2973] = 64'h801d82be01470076;
        dcache[2974] = 64'h831202eb80370000;
        dcache[2975] = 64'h017f010700530109;
        dcache[2976] = 64'h802c004f00428261;
        dcache[2977] = 64'h809c8183013c00a5;
        dcache[2978] = 64'h825c039f80690062;
        dcache[2979] = 64'h01dc003e01150150;
        dcache[2980] = 64'h806e005200d0820a;
        dcache[2981] = 64'h809e8158009f80d5;
        dcache[2982] = 64'h81bc031d00710035;
        dcache[2983] = 64'h01c50052014f00a5;
        dcache[2984] = 64'h804f00de000a81ce;
        dcache[2985] = 64'h80ef81ff00488127;
        dcache[2986] = 64'h80dc02d2015e804d;
        dcache[2987] = 64'h02a780bc008a0185;
        dcache[2988] = 64'h00350111818a0023;
        dcache[2989] = 64'h819e81be00ce81b8;
        dcache[2990] = 64'h80bd02cd01568038;
        dcache[2991] = 64'h028580b6805d0259;
        dcache[2992] = 64'h8156802d805e0088;
        dcache[2993] = 64'h801f821d00bf818f;
        dcache[2994] = 64'h804b0487005c0066;
        dcache[2995] = 64'h01a8004a01ae0133;
        dcache[2996] = 64'h8057814500ad001b;
        dcache[2997] = 64'h800a8253002d80e1;
        dcache[2998] = 64'h813e03b6803d8047;
        dcache[2999] = 64'h01e6802e005a0091;
        dcache[3000] = 64'h803780c1011b0153;
        dcache[3001] = 64'h80f2825c800d8084;
        dcache[3002] = 64'h811102f08003810e;
        dcache[3003] = 64'h024680600067014a;
        dcache[3004] = 64'h812400c6014b0129;
        dcache[3005] = 64'h006a806d0165805d;
        dcache[3006] = 64'h0028010e806c0076;
        dcache[3007] = 64'h0085002500b20185;
        dcache[3008] = 64'h811980a600878029;
        dcache[3009] = 64'h80c1811500f20034;
        dcache[3010] = 64'h80ca007480c78038;
        dcache[3011] = 64'h00748008013f0049;
        dcache[3012] = 64'h0079006880ad0014;
        dcache[3013] = 64'h8027803580c5008e;
        dcache[3014] = 64'h80838001002e8049;
        dcache[3015] = 64'h0015008080c30035;
        dcache[3016] = 64'h8013801f00468046;
        dcache[3017] = 64'h002a004580328014;
        dcache[3018] = 64'h8058001c002c801d;
        dcache[3019] = 64'h00178042802d8033;
        dcache[3020] = 64'h00050001802f0026;
        dcache[3021] = 64'h80040011803c0053;
        dcache[3022] = 64'h8027804b00128024;
        dcache[3023] = 64'h803f8046000a8041;
        dcache[3024] = 64'h002400398031804c;
        dcache[3025] = 64'h0035002f00580057;
        dcache[3026] = 64'h8046802e80200017;
        dcache[3027] = 64'h0014005200580035;
        dcache[3028] = 64'h803a802380550005;
        dcache[3029] = 64'h0003804f80058051;
        dcache[3030] = 64'h800e80260020803f;
        dcache[3031] = 64'h004780388016802f;
        dcache[3032] = 64'h803b804380008007;
        dcache[3033] = 64'h804500110041802a;
        dcache[3034] = 64'h80078037800c0054;
        dcache[3035] = 64'h003100148004803f;
        dcache[3036] = 64'h800f800480220020;
        dcache[3037] = 64'h80240026000d0014;
        dcache[3038] = 64'h80128041000a000f;
        dcache[3039] = 64'h8041001d8016801b;
        dcache[3040] = 64'h00a100538124000c;
        dcache[3041] = 64'h80a400188066006d;
        dcache[3042] = 64'h808580a800f9805c;
        dcache[3043] = 64'h00a900df80e0004f;
        dcache[3044] = 64'h01c901ad81348016;
        dcache[3045] = 64'h80de800f8167001a;
        dcache[3046] = 64'h8129815501c58121;
        dcache[3047] = 64'h013d015381898006;
        dcache[3048] = 64'h8062803881be8047;
        dcache[3049] = 64'h8015813a00bc002b;
        dcache[3050] = 64'h806d003d01700008;
        dcache[3051] = 64'h0195806e0064000b;
        dcache[3052] = 64'h80f9801a81a18050;
        dcache[3053] = 64'h800c815500c4005a;
        dcache[3054] = 64'h0037007a012e0005;
        dcache[3055] = 64'h01ad803c00cd0061;
        dcache[3056] = 64'h80a3803e819e8059;
        dcache[3057] = 64'h001b80f7010300c1;
        dcache[3058] = 64'h8024012a00f08004;
        dcache[3059] = 64'h0150806e0092803f;
        dcache[3060] = 64'h805c807800a4802d;
        dcache[3061] = 64'h007081de00fe017d;
        dcache[3062] = 64'h000401640131801f;
        dcache[3063] = 64'h01698095003e8121;
        dcache[3064] = 64'h0094006c80468116;
        dcache[3065] = 64'h8084825000d201b6;
        dcache[3066] = 64'h811a019c01bc8142;
        dcache[3067] = 64'h018880af00730141;
        dcache[3068] = 64'h80a1806100b58124;
        dcache[3069] = 64'h001e819e00af0306;
        dcache[3070] = 64'h0020024100ad0065;
        dcache[3071] = 64'h00f300ae011f010b;
        dcache[3072] = 64'h814c80f0008a8119;
        dcache[3073] = 64'h00a9828f015802c0;
        dcache[3074] = 64'h00f601d1803a00fd;
        dcache[3075] = 64'h00f90034014c00ea;
        dcache[3076] = 64'h0225021181a781b5;
        dcache[3077] = 64'h80bc81e4803e036f;
        dcache[3078] = 64'h80ea007c02be820e;
        dcache[3079] = 64'h02a1000b81380147;
        dcache[3080] = 64'h80aa004901af81bc;
        dcache[3081] = 64'h80e082d9026b02aa;
        dcache[3082] = 64'h816d02b002bb81ea;
        dcache[3083] = 64'h0382820e000e0090;
        dcache[3084] = 64'h80c980de01598227;
        dcache[3085] = 64'h008281e501c702da;
        dcache[3086] = 64'h814c01fc00968078;
        dcache[3087] = 64'h0168800a00ce0026;
        dcache[3088] = 64'h0000807500da8241;
        dcache[3089] = 64'h015a809a0118021e;
        dcache[3090] = 64'h8014023800740005;
        dcache[3091] = 64'h013c801080068006;
        dcache[3092] = 64'h00d900f180608232;
        dcache[3093] = 64'h00d881ab012a0110;
        dcache[3094] = 64'h804c01760257809d;
        dcache[3095] = 64'h030680b18116008c;
        dcache[3096] = 64'h005280458035818f;
        dcache[3097] = 64'h011181b900db8077;
        dcache[3098] = 64'h811c0117013b005c;
        dcache[3099] = 64'h025c8099802b0017;
        dcache[3100] = 64'h0087001c80768184;
        dcache[3101] = 64'h00fa814501558048;
        dcache[3102] = 64'h804800930191807e;
        dcache[3103] = 64'h02438090000c806e;
        dcache[3104] = 64'h8011811d0132810b;
        dcache[3105] = 64'h017e804f00d1804a;
        dcache[3106] = 64'h012a018280548122;
        dcache[3107] = 64'h0144807e005b801f;
        dcache[3108] = 64'h0097814f01d980c4;
        dcache[3109] = 64'h806b803380c0806a;
        dcache[3110] = 64'h810e014600188150;
        dcache[3111] = 64'h017680f180de8061;
        dcache[3112] = 64'h00b58116016c809e;
        dcache[3113] = 64'h80488035811e80eb;
        dcache[3114] = 64'h80e700e78028818d;
        dcache[3115] = 64'h019480cd808a8015;
        dcache[3116] = 64'h019600a300008048;
        dcache[3117] = 64'h81a9004d80518032;
        dcache[3118] = 64'h80bf813c004680a1;
        dcache[3119] = 64'h0188007c81718024;
        dcache[3120] = 64'h802a0051804f0021;
        dcache[3121] = 64'h001d002800388045;
        dcache[3122] = 64'h8040802f8042002e;
        dcache[3123] = 64'h801b0058800c0021;
        dcache[3124] = 64'h0048802800378028;
        dcache[3125] = 64'h0040801e00578035;
        dcache[3126] = 64'h80230047801f0007;
        dcache[3127] = 64'h8013000280360043;
        dcache[3128] = 64'h002e0043004e800e;
        dcache[3129] = 64'h8048004880240050;
        dcache[3130] = 64'h804f803680340056;
        dcache[3131] = 64'h004c000f004e8027;
        dcache[3132] = 64'h0053004f001b8039;
        dcache[3133] = 64'h8057002000468027;
        dcache[3134] = 64'h802a800e00290054;
        dcache[3135] = 64'h001a002a801e004d;
        dcache[3136] = 64'h8185007f000d8380;
        dcache[3137] = 64'h027680118310036b;
        dcache[3138] = 64'h82ca80d300000000;
        dcache[3139] = 64'h838181ec016f0267;
        dcache[3140] = 64'h80890255849c010a;
        dcache[3141] = 64'h00ad82c900000000;
        dcache[3142] = 64'h830d027b00c800e3;
        dcache[3143] = 64'h0052838283468144;
        dcache[3144] = 64'h01fc013300000000;
        dcache[3145] = 64'h002503ef00208065;
        dcache[3146] = 64'h856a036c01778228;
        dcache[3147] = 64'h82c5820e00000000;
        dcache[3148] = 64'h82bf812d01bf81fc;
        dcache[3149] = 64'h02ab00af00db006d;
        dcache[3150] = 64'h0131019400000000;
        dcache[3151] = 64'h80d50156020e013b;
        dcache[3152] = 64'h0035012201f480ea;
        dcache[3153] = 64'h8092864e00000000;
        dcache[3154] = 64'h01d4824e02088182;
        dcache[3155] = 64'h006a80e400078031;
        dcache[3156] = 64'h8590024d00000000;
        dcache[3157] = 64'h847d02510274023e;
        dcache[3158] = 64'h849181c184d90325;
        dcache[3159] = 64'h83bc872600000000;
        dcache[3160] = 64'h024f832e00378355;
        dcache[3161] = 64'h00b981e601958276;
        dcache[3162] = 64'h0176808400000000;
        dcache[3163] = 64'h818d011b815e0057;
        dcache[3164] = 64'h834d00e000d7806d;
        dcache[3165] = 64'h802b00c200000000;
        dcache[3166] = 64'h01b8015b018b81c1;
        dcache[3167] = 64'h808284f401bc01e2;
        dcache[3168] = 64'h0113009400000000;
        dcache[3169] = 64'h81ee820083ba011e;
        dcache[3170] = 64'h0155803700ee818a;
        dcache[3171] = 64'h8080003700000000;
        dcache[3172] = 64'h0109845380b50047;
        dcache[3173] = 64'h825481e183ea00c1;
        dcache[3174] = 64'h825c008f00000000;
        dcache[3175] = 64'h005d0261835581bc;
        dcache[3176] = 64'h011b02a181ab0013;
        dcache[3177] = 64'h012500b900000000;
        dcache[3178] = 64'h8175834e811d01da;
        dcache[3179] = 64'h014301da827980e8;
        dcache[3180] = 64'h02c501e800000000;
        dcache[3181] = 64'h014f82290184001a;
        dcache[3182] = 64'h86e080098206811d;
        dcache[3183] = 64'h812282b000000000;
        dcache[3184] = 64'h02a1812681d70154;
        dcache[3185] = 64'h00c00103004d80c5;
        dcache[3186] = 64'h80b5013b006300de;
        dcache[3187] = 64'h803e025480b2812b;
        dcache[3188] = 64'h8110015781598193;
        dcache[3189] = 64'h0123027c004100ea;
        dcache[3190] = 64'h822d004700000000;
        dcache[3191] = 64'h0000000000000000;
    end

    initial begin
        $dumpfile("main_tb.vcd");
        $dumpvars(0, dcache[0]);
        $dumpvars(0, dcache[1]);
        $dumpvars(0, dcache[2]);
        $dumpvars(0, dcache[3]);
        $dumpvars(0, dcache[4]);
        $dumpvars(0, dcache[5]);
        $dumpvars(0, dcache[6]);
        $dumpvars(0, dcache[7]);
        $dumpvars(0, dcache[8]);
        $dumpvars(0, dcache[9]);
        $dumpvars(0, dcache[10]);
        $dumpvars(0, dcache[11]);
        $dumpvars(0, dcache[12]);
        $dumpvars(0, dcache[13]);
        $dumpvars(0, dcache[14]);
        $dumpvars(0, dcache[15]);
        $dumpvars(0, dcache[16]);
        $dumpvars(0, dcache[17]);
        $dumpvars(0, dcache[18]);
        $dumpvars(0, dcache[19]);
        $dumpvars(0, dcache[20]);
        $dumpvars(0, dcache[21]);
        $dumpvars(0, dcache[22]);
        $dumpvars(0, dcache[23]);
        $dumpvars(0, dcache[24]);
        $dumpvars(0, dcache[25]);
        $dumpvars(0, dcache[26]);
        $dumpvars(0, dcache[27]);
        $dumpvars(0, dcache[28]);
        $dumpvars(0, dcache[29]);
        $dumpvars(0, dcache[30]);
        $dumpvars(0, dcache[31]);
        $dumpvars(0, dcache[32]);
        $dumpvars(0, dcache[33]);
        $dumpvars(0, dcache[34]);
        $dumpvars(0, dcache[35]);
        $dumpvars(0, dcache[36]);
        $dumpvars(0, dcache[37]);
        $dumpvars(0, dcache[38]);
        $dumpvars(0, dcache[39]);
        $dumpvars(0, dcache[40]);
        $dumpvars(0, dcache[41]);
        $dumpvars(0, dcache[42]);
        $dumpvars(0, dcache[43]);
        $dumpvars(0, dcache[44]);
        $dumpvars(0, dcache[45]);
        $dumpvars(0, dcache[46]);
        $dumpvars(0, dcache[47]);
        $dumpvars(0, dcache[48]);
        $dumpvars(0, dcache[49]);
        $dumpvars(0, dcache[50]);
        $dumpvars(0, dcache[51]);
        $dumpvars(0, dcache[52]);
        $dumpvars(0, dcache[53]);
        $dumpvars(0, dcache[54]);
        $dumpvars(0, dcache[55]);
        $dumpvars(0, dcache[56]);
        $dumpvars(0, dcache[57]);
        $dumpvars(0, dcache[58]);
        $dumpvars(0, dcache[59]);
        $dumpvars(0, dcache[60]);
        $dumpvars(0, dcache[61]);
        $dumpvars(0, dcache[62]);
        $dumpvars(0, dcache[63]);
        $dumpvars(0, dcache[64]);
        $dumpvars(0, dcache[65]);
        $dumpvars(0, dcache[66]);
        $dumpvars(0, dcache[67]);
        $dumpvars(0, dcache[68]);
        $dumpvars(0, dcache[69]);
        $dumpvars(0, dcache[70]);
        $dumpvars(0, dcache[71]);
        $dumpvars(0, dcache[72]);
        $dumpvars(0, dcache[73]);
        $dumpvars(0, dcache[74]);
        $dumpvars(0, dcache[75]);
        $dumpvars(0, dcache[76]);
        $dumpvars(0, dcache[77]);
        $dumpvars(0, dcache[78]);
        $dumpvars(0, dcache[79]);
        $dumpvars(0, dcache[80]);
        $dumpvars(0, dcache[81]);
        $dumpvars(0, dcache[82]);
        $dumpvars(0, dcache[83]);
        $dumpvars(0, dcache[84]);
        $dumpvars(0, dcache[85]);
        $dumpvars(0, dcache[86]);
        $dumpvars(0, dcache[87]);
        $dumpvars(0, dcache[88]);
        $dumpvars(0, dcache[89]);
        $dumpvars(0, dcache[90]);
        $dumpvars(0, dcache[91]);
        $dumpvars(0, dcache[92]);
        $dumpvars(0, dcache[93]);
        $dumpvars(0, dcache[94]);
        $dumpvars(0, dcache[95]);
        $dumpvars(0, dcache[96]);
        $dumpvars(0, dcache[97]);
        $dumpvars(0, dcache[98]);
        $dumpvars(0, dcache[99]);
        $dumpvars(0, dcache[100]);
        $dumpvars(0, dcache[101]);
        $dumpvars(0, dcache[102]);
        $dumpvars(0, dcache[103]);
        $dumpvars(0, dcache[104]);
        $dumpvars(0, dcache[105]);
        $dumpvars(0, dcache[106]);
        $dumpvars(0, dcache[107]);
        $dumpvars(0, dcache[108]);
        $dumpvars(0, dcache[109]);
        $dumpvars(0, dcache[110]);
        $dumpvars(0, dcache[111]);
        $dumpvars(0, dcache[112]);
        $dumpvars(0, dcache[113]);
        $dumpvars(0, dcache[114]);
        $dumpvars(0, dcache[115]);
        $dumpvars(0, dcache[116]);
        $dumpvars(0, dcache[117]);
        $dumpvars(0, dcache[118]);
        $dumpvars(0, dcache[119]);
        $dumpvars(0, dcache[120]);
        $dumpvars(0, dcache[121]);
        $dumpvars(0, dcache[122]);
        $dumpvars(0, dcache[123]);
        $dumpvars(0, dcache[124]);
        $dumpvars(0, dcache[125]);
        $dumpvars(0, dcache[126]);
        $dumpvars(0, dcache[127]);
    end

endmodule
